VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_rejunity_z80
  CLASS BLOCK ;
  FOREIGN tt_um_rejunity_z80 ;
  ORIGIN 0.000 0.000 ;
  SIZE 711.200 BY 325.360 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 3.620 23.780 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 61.050 3.620 62.650 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.920 3.620 101.520 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.790 3.620 140.390 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 177.660 3.620 179.260 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 216.530 3.620 218.130 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 255.400 3.620 257.000 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 294.270 3.620 295.870 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 333.140 3.620 334.740 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 372.010 3.620 373.610 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 410.880 3.620 412.480 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.750 3.620 451.350 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 488.620 3.620 490.220 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 527.490 3.620 529.090 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 566.360 3.620 567.960 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.230 3.620 606.830 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 644.100 3.620 645.700 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 682.970 3.620 684.570 321.740 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 3.620 20.480 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 57.750 3.620 59.350 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 96.620 3.620 98.220 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 135.490 3.620 137.090 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 174.360 3.620 175.960 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 213.230 3.620 214.830 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.100 3.620 253.700 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 290.970 3.620 292.570 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.840 3.620 331.440 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 368.710 3.620 370.310 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 407.580 3.620 409.180 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 446.450 3.620 448.050 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 485.320 3.620 486.920 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 524.190 3.620 525.790 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 563.060 3.620 564.660 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 601.930 3.620 603.530 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 640.800 3.620 642.400 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 679.670 3.620 681.270 321.740 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    PORT
      LAYER Metal4 ;
        RECT 331.090 324.360 331.390 325.360 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal4 ;
        RECT 338.370 324.360 338.670 325.360 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 323.810 324.360 324.110 325.360 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 316.530 324.360 316.830 325.360 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    PORT
      LAYER Metal4 ;
        RECT 309.250 324.360 309.550 325.360 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    PORT
      LAYER Metal4 ;
        RECT 301.970 324.360 302.270 325.360 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 294.690 324.360 294.990 325.360 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    PORT
      LAYER Metal4 ;
        RECT 287.410 324.360 287.710 325.360 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 280.130 324.360 280.430 325.360 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    PORT
      LAYER Metal4 ;
        RECT 272.850 324.360 273.150 325.360 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    PORT
      LAYER Metal4 ;
        RECT 265.570 324.360 265.870 325.360 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 258.290 324.360 258.590 325.360 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 251.010 324.360 251.310 325.360 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 243.730 324.360 244.030 325.360 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 236.450 324.360 236.750 325.360 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 229.170 324.360 229.470 325.360 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 221.890 324.360 222.190 325.360 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 214.610 324.360 214.910 325.360 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 207.330 324.360 207.630 325.360 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal4 ;
        RECT 83.570 324.360 83.870 325.360 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal4 ;
        RECT 76.290 324.360 76.590 325.360 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal4 ;
        RECT 69.010 324.360 69.310 325.360 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal4 ;
        RECT 61.730 324.360 62.030 325.360 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal4 ;
        RECT 54.450 324.360 54.750 325.360 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal4 ;
        RECT 47.170 324.360 47.470 325.360 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal4 ;
        RECT 39.890 324.360 40.190 325.360 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal4 ;
        RECT 32.610 324.360 32.910 325.360 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.114000 ;
    ANTENNADIFFAREA 2.111200 ;
    PORT
      LAYER Metal4 ;
        RECT 141.810 324.360 142.110 325.360 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.114000 ;
    ANTENNADIFFAREA 2.111200 ;
    PORT
      LAYER Metal4 ;
        RECT 134.530 324.360 134.830 325.360 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.114000 ;
    ANTENNADIFFAREA 2.111200 ;
    PORT
      LAYER Metal4 ;
        RECT 127.250 324.360 127.550 325.360 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.199000 ;
    ANTENNADIFFAREA 2.111200 ;
    PORT
      LAYER Metal4 ;
        RECT 119.970 324.360 120.270 325.360 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal4 ;
        RECT 112.690 324.360 112.990 325.360 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.199000 ;
    ANTENNADIFFAREA 2.111200 ;
    PORT
      LAYER Metal4 ;
        RECT 105.410 324.360 105.710 325.360 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.133000 ;
    ANTENNADIFFAREA 2.111200 ;
    PORT
      LAYER Metal4 ;
        RECT 98.130 324.360 98.430 325.360 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898000 ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal4 ;
        RECT 90.850 324.360 91.150 325.360 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.030500 ;
    PORT
      LAYER Metal4 ;
        RECT 200.050 324.360 200.350 325.360 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.369000 ;
    PORT
      LAYER Metal4 ;
        RECT 192.770 324.360 193.070 325.360 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.030500 ;
    PORT
      LAYER Metal4 ;
        RECT 185.490 324.360 185.790 325.360 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.389000 ;
    PORT
      LAYER Metal4 ;
        RECT 178.210 324.360 178.510 325.360 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.369000 ;
    PORT
      LAYER Metal4 ;
        RECT 170.930 324.360 171.230 325.360 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.369000 ;
    PORT
      LAYER Metal4 ;
        RECT 163.650 324.360 163.950 325.360 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.369000 ;
    PORT
      LAYER Metal4 ;
        RECT 156.370 324.360 156.670 325.360 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.369000 ;
    PORT
      LAYER Metal4 ;
        RECT 149.090 324.360 149.390 325.360 ;
    END
  END uo_out[7]
  OBS
      LAYER Nwell ;
        RECT 2.930 319.280 708.270 321.870 ;
      LAYER Pwell ;
        RECT 2.930 315.760 708.270 319.280 ;
      LAYER Nwell ;
        RECT 2.930 311.440 708.270 315.760 ;
      LAYER Pwell ;
        RECT 2.930 307.920 708.270 311.440 ;
      LAYER Nwell ;
        RECT 2.930 303.600 708.270 307.920 ;
      LAYER Pwell ;
        RECT 2.930 300.080 708.270 303.600 ;
      LAYER Nwell ;
        RECT 2.930 295.760 708.270 300.080 ;
      LAYER Pwell ;
        RECT 2.930 292.240 708.270 295.760 ;
      LAYER Nwell ;
        RECT 2.930 287.920 708.270 292.240 ;
      LAYER Pwell ;
        RECT 2.930 284.400 708.270 287.920 ;
      LAYER Nwell ;
        RECT 2.930 280.080 708.270 284.400 ;
      LAYER Pwell ;
        RECT 2.930 276.560 708.270 280.080 ;
      LAYER Nwell ;
        RECT 2.930 272.240 708.270 276.560 ;
      LAYER Pwell ;
        RECT 2.930 268.720 708.270 272.240 ;
      LAYER Nwell ;
        RECT 2.930 264.400 708.270 268.720 ;
      LAYER Pwell ;
        RECT 2.930 260.880 708.270 264.400 ;
      LAYER Nwell ;
        RECT 2.930 256.560 708.270 260.880 ;
      LAYER Pwell ;
        RECT 2.930 253.040 708.270 256.560 ;
      LAYER Nwell ;
        RECT 2.930 248.720 708.270 253.040 ;
      LAYER Pwell ;
        RECT 2.930 245.200 708.270 248.720 ;
      LAYER Nwell ;
        RECT 2.930 240.880 708.270 245.200 ;
      LAYER Pwell ;
        RECT 2.930 237.360 708.270 240.880 ;
      LAYER Nwell ;
        RECT 2.930 233.040 708.270 237.360 ;
      LAYER Pwell ;
        RECT 2.930 229.520 708.270 233.040 ;
      LAYER Nwell ;
        RECT 2.930 225.200 708.270 229.520 ;
      LAYER Pwell ;
        RECT 2.930 221.680 708.270 225.200 ;
      LAYER Nwell ;
        RECT 2.930 217.360 708.270 221.680 ;
      LAYER Pwell ;
        RECT 2.930 213.840 708.270 217.360 ;
      LAYER Nwell ;
        RECT 2.930 209.520 708.270 213.840 ;
      LAYER Pwell ;
        RECT 2.930 206.000 708.270 209.520 ;
      LAYER Nwell ;
        RECT 2.930 201.680 708.270 206.000 ;
      LAYER Pwell ;
        RECT 2.930 198.160 708.270 201.680 ;
      LAYER Nwell ;
        RECT 2.930 193.840 708.270 198.160 ;
      LAYER Pwell ;
        RECT 2.930 190.320 708.270 193.840 ;
      LAYER Nwell ;
        RECT 2.930 186.000 708.270 190.320 ;
      LAYER Pwell ;
        RECT 2.930 182.480 708.270 186.000 ;
      LAYER Nwell ;
        RECT 2.930 178.160 708.270 182.480 ;
      LAYER Pwell ;
        RECT 2.930 174.640 708.270 178.160 ;
      LAYER Nwell ;
        RECT 2.930 170.320 708.270 174.640 ;
      LAYER Pwell ;
        RECT 2.930 166.800 708.270 170.320 ;
      LAYER Nwell ;
        RECT 2.930 162.480 708.270 166.800 ;
      LAYER Pwell ;
        RECT 2.930 158.960 708.270 162.480 ;
      LAYER Nwell ;
        RECT 2.930 154.640 708.270 158.960 ;
      LAYER Pwell ;
        RECT 2.930 151.120 708.270 154.640 ;
      LAYER Nwell ;
        RECT 2.930 146.800 708.270 151.120 ;
      LAYER Pwell ;
        RECT 2.930 143.280 708.270 146.800 ;
      LAYER Nwell ;
        RECT 2.930 138.960 708.270 143.280 ;
      LAYER Pwell ;
        RECT 2.930 135.440 708.270 138.960 ;
      LAYER Nwell ;
        RECT 2.930 131.120 708.270 135.440 ;
      LAYER Pwell ;
        RECT 2.930 127.600 708.270 131.120 ;
      LAYER Nwell ;
        RECT 2.930 123.280 708.270 127.600 ;
      LAYER Pwell ;
        RECT 2.930 119.760 708.270 123.280 ;
      LAYER Nwell ;
        RECT 2.930 115.440 708.270 119.760 ;
      LAYER Pwell ;
        RECT 2.930 111.920 708.270 115.440 ;
      LAYER Nwell ;
        RECT 2.930 107.600 708.270 111.920 ;
      LAYER Pwell ;
        RECT 2.930 104.080 708.270 107.600 ;
      LAYER Nwell ;
        RECT 2.930 99.760 708.270 104.080 ;
      LAYER Pwell ;
        RECT 2.930 96.240 708.270 99.760 ;
      LAYER Nwell ;
        RECT 2.930 91.920 708.270 96.240 ;
      LAYER Pwell ;
        RECT 2.930 88.400 708.270 91.920 ;
      LAYER Nwell ;
        RECT 2.930 84.080 708.270 88.400 ;
      LAYER Pwell ;
        RECT 2.930 80.560 708.270 84.080 ;
      LAYER Nwell ;
        RECT 2.930 76.240 708.270 80.560 ;
      LAYER Pwell ;
        RECT 2.930 72.720 708.270 76.240 ;
      LAYER Nwell ;
        RECT 2.930 68.400 708.270 72.720 ;
      LAYER Pwell ;
        RECT 2.930 64.880 708.270 68.400 ;
      LAYER Nwell ;
        RECT 2.930 60.560 708.270 64.880 ;
      LAYER Pwell ;
        RECT 2.930 57.040 708.270 60.560 ;
      LAYER Nwell ;
        RECT 2.930 52.720 708.270 57.040 ;
      LAYER Pwell ;
        RECT 2.930 49.200 708.270 52.720 ;
      LAYER Nwell ;
        RECT 2.930 44.880 708.270 49.200 ;
      LAYER Pwell ;
        RECT 2.930 41.360 708.270 44.880 ;
      LAYER Nwell ;
        RECT 2.930 37.040 708.270 41.360 ;
      LAYER Pwell ;
        RECT 2.930 33.520 708.270 37.040 ;
      LAYER Nwell ;
        RECT 2.930 29.200 708.270 33.520 ;
      LAYER Pwell ;
        RECT 2.930 25.680 708.270 29.200 ;
      LAYER Nwell ;
        RECT 2.930 21.360 708.270 25.680 ;
      LAYER Pwell ;
        RECT 2.930 17.840 708.270 21.360 ;
      LAYER Nwell ;
        RECT 2.930 13.520 708.270 17.840 ;
      LAYER Pwell ;
        RECT 2.930 10.000 708.270 13.520 ;
      LAYER Nwell ;
        RECT 2.930 5.680 708.270 10.000 ;
      LAYER Pwell ;
        RECT 2.930 3.490 708.270 5.680 ;
      LAYER Metal1 ;
        RECT 3.360 3.620 707.840 321.740 ;
      LAYER Metal2 ;
        RECT 3.500 0.090 697.620 324.710 ;
      LAYER Metal3 ;
        RECT 3.450 0.140 697.670 325.220 ;
      LAYER Metal4 ;
        RECT 9.660 324.060 32.310 325.270 ;
        RECT 33.210 324.060 39.590 325.270 ;
        RECT 40.490 324.060 46.870 325.270 ;
        RECT 47.770 324.060 54.150 325.270 ;
        RECT 55.050 324.060 61.430 325.270 ;
        RECT 62.330 324.060 68.710 325.270 ;
        RECT 69.610 324.060 75.990 325.270 ;
        RECT 76.890 324.060 83.270 325.270 ;
        RECT 84.170 324.060 90.550 325.270 ;
        RECT 91.450 324.060 97.830 325.270 ;
        RECT 98.730 324.060 105.110 325.270 ;
        RECT 106.010 324.060 112.390 325.270 ;
        RECT 113.290 324.060 119.670 325.270 ;
        RECT 120.570 324.060 126.950 325.270 ;
        RECT 127.850 324.060 134.230 325.270 ;
        RECT 135.130 324.060 141.510 325.270 ;
        RECT 142.410 324.060 148.790 325.270 ;
        RECT 149.690 324.060 156.070 325.270 ;
        RECT 156.970 324.060 163.350 325.270 ;
        RECT 164.250 324.060 170.630 325.270 ;
        RECT 171.530 324.060 177.910 325.270 ;
        RECT 178.810 324.060 185.190 325.270 ;
        RECT 186.090 324.060 192.470 325.270 ;
        RECT 193.370 324.060 199.750 325.270 ;
        RECT 200.650 324.060 207.030 325.270 ;
        RECT 207.930 324.060 214.310 325.270 ;
        RECT 215.210 324.060 221.590 325.270 ;
        RECT 222.490 324.060 228.870 325.270 ;
        RECT 229.770 324.060 236.150 325.270 ;
        RECT 237.050 324.060 243.430 325.270 ;
        RECT 244.330 324.060 250.710 325.270 ;
        RECT 251.610 324.060 257.990 325.270 ;
        RECT 258.890 324.060 265.270 325.270 ;
        RECT 266.170 324.060 272.550 325.270 ;
        RECT 273.450 324.060 279.830 325.270 ;
        RECT 280.730 324.060 287.110 325.270 ;
        RECT 288.010 324.060 294.390 325.270 ;
        RECT 295.290 324.060 301.670 325.270 ;
        RECT 302.570 324.060 308.950 325.270 ;
        RECT 309.850 324.060 316.230 325.270 ;
        RECT 317.130 324.060 323.510 325.270 ;
        RECT 324.410 324.060 330.790 325.270 ;
        RECT 331.690 324.060 338.070 325.270 ;
        RECT 338.970 324.060 662.900 325.270 ;
        RECT 9.660 322.040 662.900 324.060 ;
        RECT 9.660 3.320 18.580 322.040 ;
        RECT 20.780 3.320 21.880 322.040 ;
        RECT 24.080 3.320 57.450 322.040 ;
        RECT 59.650 3.320 60.750 322.040 ;
        RECT 62.950 3.320 96.320 322.040 ;
        RECT 98.520 3.320 99.620 322.040 ;
        RECT 101.820 3.320 135.190 322.040 ;
        RECT 137.390 3.320 138.490 322.040 ;
        RECT 140.690 3.320 174.060 322.040 ;
        RECT 176.260 3.320 177.360 322.040 ;
        RECT 179.560 3.320 212.930 322.040 ;
        RECT 215.130 3.320 216.230 322.040 ;
        RECT 218.430 3.320 251.800 322.040 ;
        RECT 254.000 3.320 255.100 322.040 ;
        RECT 257.300 3.320 290.670 322.040 ;
        RECT 292.870 3.320 293.970 322.040 ;
        RECT 296.170 3.320 329.540 322.040 ;
        RECT 331.740 3.320 332.840 322.040 ;
        RECT 335.040 3.320 368.410 322.040 ;
        RECT 370.610 3.320 371.710 322.040 ;
        RECT 373.910 3.320 407.280 322.040 ;
        RECT 409.480 3.320 410.580 322.040 ;
        RECT 412.780 3.320 446.150 322.040 ;
        RECT 448.350 3.320 449.450 322.040 ;
        RECT 451.650 3.320 485.020 322.040 ;
        RECT 487.220 3.320 488.320 322.040 ;
        RECT 490.520 3.320 523.890 322.040 ;
        RECT 526.090 3.320 527.190 322.040 ;
        RECT 529.390 3.320 562.760 322.040 ;
        RECT 564.960 3.320 566.060 322.040 ;
        RECT 568.260 3.320 601.630 322.040 ;
        RECT 603.830 3.320 604.930 322.040 ;
        RECT 607.130 3.320 640.500 322.040 ;
        RECT 642.700 3.320 643.800 322.040 ;
        RECT 646.000 3.320 662.900 322.040 ;
        RECT 9.660 0.090 662.900 3.320 ;
  END
END tt_um_rejunity_z80
END LIBRARY

