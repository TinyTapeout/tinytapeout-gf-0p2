VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_urish_simon
  CLASS BLOCK ;
  FOREIGN tt_um_urish_simon ;
  ORIGIN 0.000 0.000 ;
  SIZE 346.640 BY 160.720 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 3.620 23.780 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 61.050 3.620 62.650 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.920 3.620 101.520 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.790 3.620 140.390 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 177.660 3.620 179.260 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 216.530 3.620 218.130 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 255.400 3.620 257.000 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 294.270 3.620 295.870 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 333.140 3.620 334.740 157.100 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 3.620 20.480 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 57.750 3.620 59.350 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 96.620 3.620 98.220 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 135.490 3.620 137.090 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 174.360 3.620 175.960 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 213.230 3.620 214.830 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.100 3.620 253.700 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 290.970 3.620 292.570 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.840 3.620 331.440 157.100 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 330.810 159.720 331.110 160.720 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 338.090 159.720 338.390 160.720 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 323.530 159.720 323.830 160.720 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 316.250 159.720 316.550 160.720 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    PORT
      LAYER Metal4 ;
        RECT 308.970 159.720 309.270 160.720 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 301.690 159.720 301.990 160.720 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    PORT
      LAYER Metal4 ;
        RECT 294.410 159.720 294.710 160.720 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    PORT
      LAYER Metal4 ;
        RECT 287.130 159.720 287.430 160.720 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 279.850 159.720 280.150 160.720 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 272.570 159.720 272.870 160.720 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 265.290 159.720 265.590 160.720 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 258.010 159.720 258.310 160.720 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 250.730 159.720 251.030 160.720 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 243.450 159.720 243.750 160.720 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 236.170 159.720 236.470 160.720 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 228.890 159.720 229.190 160.720 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 221.610 159.720 221.910 160.720 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 214.330 159.720 214.630 160.720 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 207.050 159.720 207.350 160.720 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal4 ;
        RECT 83.290 159.720 83.590 160.720 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal4 ;
        RECT 76.010 159.720 76.310 160.720 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal4 ;
        RECT 68.730 159.720 69.030 160.720 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal4 ;
        RECT 61.450 159.720 61.750 160.720 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal4 ;
        RECT 54.170 159.720 54.470 160.720 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal4 ;
        RECT 46.890 159.720 47.190 160.720 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal4 ;
        RECT 39.610 159.720 39.910 160.720 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 32.330 159.720 32.630 160.720 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal4 ;
        RECT 141.530 159.720 141.830 160.720 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal4 ;
        RECT 134.250 159.720 134.550 160.720 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal4 ;
        RECT 126.970 159.720 127.270 160.720 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal4 ;
        RECT 119.690 159.720 119.990 160.720 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal4 ;
        RECT 112.410 159.720 112.710 160.720 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal4 ;
        RECT 105.130 159.720 105.430 160.720 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal4 ;
        RECT 97.850 159.720 98.150 160.720 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 90.570 159.720 90.870 160.720 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal4 ;
        RECT 199.770 159.720 200.070 160.720 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal4 ;
        RECT 192.490 159.720 192.790 160.720 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal4 ;
        RECT 185.210 159.720 185.510 160.720 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal4 ;
        RECT 177.930 159.720 178.230 160.720 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal4 ;
        RECT 170.650 159.720 170.950 160.720 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal4 ;
        RECT 163.370 159.720 163.670 160.720 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.060800 ;
    PORT
      LAYER Metal4 ;
        RECT 156.090 159.720 156.390 160.720 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal4 ;
        RECT 148.810 159.720 149.110 160.720 ;
    END
  END uo_out[7]
  OBS
      LAYER Nwell ;
        RECT 2.930 154.640 343.710 157.230 ;
      LAYER Pwell ;
        RECT 2.930 151.120 343.710 154.640 ;
      LAYER Nwell ;
        RECT 2.930 146.800 343.710 151.120 ;
      LAYER Pwell ;
        RECT 2.930 143.280 343.710 146.800 ;
      LAYER Nwell ;
        RECT 2.930 138.960 343.710 143.280 ;
      LAYER Pwell ;
        RECT 2.930 135.440 343.710 138.960 ;
      LAYER Nwell ;
        RECT 2.930 131.120 343.710 135.440 ;
      LAYER Pwell ;
        RECT 2.930 127.600 343.710 131.120 ;
      LAYER Nwell ;
        RECT 2.930 123.280 343.710 127.600 ;
      LAYER Pwell ;
        RECT 2.930 119.760 343.710 123.280 ;
      LAYER Nwell ;
        RECT 2.930 115.440 343.710 119.760 ;
      LAYER Pwell ;
        RECT 2.930 111.920 343.710 115.440 ;
      LAYER Nwell ;
        RECT 2.930 107.600 343.710 111.920 ;
      LAYER Pwell ;
        RECT 2.930 104.080 343.710 107.600 ;
      LAYER Nwell ;
        RECT 2.930 99.760 343.710 104.080 ;
      LAYER Pwell ;
        RECT 2.930 96.240 343.710 99.760 ;
      LAYER Nwell ;
        RECT 2.930 91.920 343.710 96.240 ;
      LAYER Pwell ;
        RECT 2.930 88.400 343.710 91.920 ;
      LAYER Nwell ;
        RECT 2.930 84.080 343.710 88.400 ;
      LAYER Pwell ;
        RECT 2.930 80.560 343.710 84.080 ;
      LAYER Nwell ;
        RECT 2.930 76.240 343.710 80.560 ;
      LAYER Pwell ;
        RECT 2.930 72.720 343.710 76.240 ;
      LAYER Nwell ;
        RECT 2.930 68.400 343.710 72.720 ;
      LAYER Pwell ;
        RECT 2.930 64.880 343.710 68.400 ;
      LAYER Nwell ;
        RECT 2.930 60.560 343.710 64.880 ;
      LAYER Pwell ;
        RECT 2.930 57.040 343.710 60.560 ;
      LAYER Nwell ;
        RECT 2.930 52.720 343.710 57.040 ;
      LAYER Pwell ;
        RECT 2.930 49.200 343.710 52.720 ;
      LAYER Nwell ;
        RECT 2.930 44.880 343.710 49.200 ;
      LAYER Pwell ;
        RECT 2.930 41.360 343.710 44.880 ;
      LAYER Nwell ;
        RECT 2.930 37.040 343.710 41.360 ;
      LAYER Pwell ;
        RECT 2.930 33.520 343.710 37.040 ;
      LAYER Nwell ;
        RECT 2.930 29.200 343.710 33.520 ;
      LAYER Pwell ;
        RECT 2.930 25.680 343.710 29.200 ;
      LAYER Nwell ;
        RECT 2.930 21.360 343.710 25.680 ;
      LAYER Pwell ;
        RECT 2.930 17.840 343.710 21.360 ;
      LAYER Nwell ;
        RECT 2.930 13.520 343.710 17.840 ;
      LAYER Pwell ;
        RECT 2.930 10.000 343.710 13.520 ;
      LAYER Nwell ;
        RECT 2.930 5.680 343.710 10.000 ;
      LAYER Pwell ;
        RECT 2.930 3.490 343.710 5.680 ;
      LAYER Metal1 ;
        RECT 3.360 3.620 343.280 157.100 ;
      LAYER Metal2 ;
        RECT 19.020 2.330 346.500 160.630 ;
      LAYER Metal3 ;
        RECT 18.970 1.820 346.550 160.580 ;
      LAYER Metal4 ;
        RECT 32.930 159.420 39.310 159.890 ;
        RECT 40.210 159.420 46.590 159.890 ;
        RECT 47.490 159.420 53.870 159.890 ;
        RECT 54.770 159.420 61.150 159.890 ;
        RECT 62.050 159.420 68.430 159.890 ;
        RECT 69.330 159.420 75.710 159.890 ;
        RECT 76.610 159.420 82.990 159.890 ;
        RECT 83.890 159.420 90.270 159.890 ;
        RECT 91.170 159.420 97.550 159.890 ;
        RECT 98.450 159.420 104.830 159.890 ;
        RECT 105.730 159.420 112.110 159.890 ;
        RECT 113.010 159.420 119.390 159.890 ;
        RECT 120.290 159.420 126.670 159.890 ;
        RECT 127.570 159.420 133.950 159.890 ;
        RECT 134.850 159.420 141.230 159.890 ;
        RECT 142.130 159.420 148.510 159.890 ;
        RECT 149.410 159.420 155.790 159.890 ;
        RECT 156.690 159.420 163.070 159.890 ;
        RECT 163.970 159.420 170.350 159.890 ;
        RECT 171.250 159.420 177.630 159.890 ;
        RECT 178.530 159.420 184.910 159.890 ;
        RECT 185.810 159.420 192.190 159.890 ;
        RECT 193.090 159.420 199.470 159.890 ;
        RECT 200.370 159.420 206.750 159.890 ;
        RECT 207.650 159.420 214.030 159.890 ;
        RECT 214.930 159.420 221.310 159.890 ;
        RECT 222.210 159.420 228.590 159.890 ;
        RECT 229.490 159.420 235.870 159.890 ;
        RECT 236.770 159.420 243.150 159.890 ;
        RECT 244.050 159.420 250.430 159.890 ;
        RECT 251.330 159.420 257.710 159.890 ;
        RECT 258.610 159.420 264.990 159.890 ;
        RECT 265.890 159.420 272.270 159.890 ;
        RECT 273.170 159.420 279.550 159.890 ;
        RECT 280.450 159.420 286.830 159.890 ;
        RECT 287.730 159.420 294.110 159.890 ;
        RECT 295.010 159.420 301.390 159.890 ;
        RECT 302.290 159.420 308.670 159.890 ;
        RECT 309.570 159.420 315.950 159.890 ;
        RECT 316.850 159.420 323.230 159.890 ;
        RECT 324.130 159.420 330.510 159.890 ;
        RECT 331.410 159.420 337.790 159.890 ;
        RECT 338.690 159.420 341.460 159.890 ;
        RECT 32.340 157.400 341.460 159.420 ;
        RECT 32.340 3.320 57.450 157.400 ;
        RECT 59.650 3.320 60.750 157.400 ;
        RECT 62.950 3.320 96.320 157.400 ;
        RECT 98.520 3.320 99.620 157.400 ;
        RECT 101.820 3.320 135.190 157.400 ;
        RECT 137.390 3.320 138.490 157.400 ;
        RECT 140.690 3.320 174.060 157.400 ;
        RECT 176.260 3.320 177.360 157.400 ;
        RECT 179.560 3.320 212.930 157.400 ;
        RECT 215.130 3.320 216.230 157.400 ;
        RECT 218.430 3.320 251.800 157.400 ;
        RECT 254.000 3.320 255.100 157.400 ;
        RECT 257.300 3.320 290.670 157.400 ;
        RECT 292.870 3.320 293.970 157.400 ;
        RECT 296.170 3.320 329.540 157.400 ;
        RECT 331.740 3.320 332.840 157.400 ;
        RECT 335.040 3.320 341.460 157.400 ;
        RECT 32.340 1.770 341.460 3.320 ;
  END
END tt_um_urish_simon
END LIBRARY

