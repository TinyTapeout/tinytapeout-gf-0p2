VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_a1k0n_nyancat
  CLASS BLOCK ;
  FOREIGN tt_um_a1k0n_nyancat ;
  ORIGIN 0.000 0.000 ;
  SIZE 346.640 BY 325.360 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 3.620 23.780 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 61.050 3.620 62.650 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.920 3.620 101.520 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.790 3.620 140.390 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 177.660 3.620 179.260 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 216.530 3.620 218.130 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 255.400 3.620 257.000 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 294.270 3.620 295.870 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 333.140 3.620 334.740 321.740 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 3.620 20.480 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 57.750 3.620 59.350 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 96.620 3.620 98.220 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 135.490 3.620 137.090 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 174.360 3.620 175.960 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 213.230 3.620 214.830 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.100 3.620 253.700 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 290.970 3.620 292.570 321.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.840 3.620 331.440 321.740 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    PORT
      LAYER Metal4 ;
        RECT 331.090 324.360 331.390 325.360 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 338.370 324.360 338.670 325.360 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    PORT
      LAYER Metal4 ;
        RECT 323.810 324.360 324.110 325.360 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 316.530 324.360 316.830 325.360 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 309.250 324.360 309.550 325.360 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 301.970 324.360 302.270 325.360 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 294.690 324.360 294.990 325.360 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 287.410 324.360 287.710 325.360 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 280.130 324.360 280.430 325.360 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 272.850 324.360 273.150 325.360 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 265.570 324.360 265.870 325.360 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 258.290 324.360 258.590 325.360 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 251.010 324.360 251.310 325.360 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 243.730 324.360 244.030 325.360 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 236.450 324.360 236.750 325.360 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 229.170 324.360 229.470 325.360 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 221.890 324.360 222.190 325.360 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 214.610 324.360 214.910 325.360 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 207.330 324.360 207.630 325.360 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 83.570 324.360 83.870 325.360 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 76.290 324.360 76.590 325.360 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 69.010 324.360 69.310 325.360 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 61.730 324.360 62.030 325.360 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 54.450 324.360 54.750 325.360 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 47.170 324.360 47.470 325.360 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 39.890 324.360 40.190 325.360 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal4 ;
        RECT 32.610 324.360 32.910 325.360 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 141.810 324.360 142.110 325.360 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 134.530 324.360 134.830 325.360 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 127.250 324.360 127.550 325.360 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 119.970 324.360 120.270 325.360 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 112.690 324.360 112.990 325.360 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 105.410 324.360 105.710 325.360 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 98.130 324.360 98.430 325.360 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 90.850 324.360 91.150 325.360 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal4 ;
        RECT 200.050 324.360 200.350 325.360 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal4 ;
        RECT 192.770 324.360 193.070 325.360 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal4 ;
        RECT 185.490 324.360 185.790 325.360 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal4 ;
        RECT 178.210 324.360 178.510 325.360 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal4 ;
        RECT 170.930 324.360 171.230 325.360 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal4 ;
        RECT 163.650 324.360 163.950 325.360 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.055600 ;
    PORT
      LAYER Metal4 ;
        RECT 156.370 324.360 156.670 325.360 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 149.090 324.360 149.390 325.360 ;
    END
  END uo_out[7]
  OBS
      LAYER Nwell ;
        RECT 2.930 319.280 343.710 321.870 ;
      LAYER Pwell ;
        RECT 2.930 315.760 343.710 319.280 ;
      LAYER Nwell ;
        RECT 2.930 311.440 343.710 315.760 ;
      LAYER Pwell ;
        RECT 2.930 307.920 343.710 311.440 ;
      LAYER Nwell ;
        RECT 2.930 303.600 343.710 307.920 ;
      LAYER Pwell ;
        RECT 2.930 300.080 343.710 303.600 ;
      LAYER Nwell ;
        RECT 2.930 295.760 343.710 300.080 ;
      LAYER Pwell ;
        RECT 2.930 292.240 343.710 295.760 ;
      LAYER Nwell ;
        RECT 2.930 287.920 343.710 292.240 ;
      LAYER Pwell ;
        RECT 2.930 284.400 343.710 287.920 ;
      LAYER Nwell ;
        RECT 2.930 280.080 343.710 284.400 ;
      LAYER Pwell ;
        RECT 2.930 276.560 343.710 280.080 ;
      LAYER Nwell ;
        RECT 2.930 272.240 343.710 276.560 ;
      LAYER Pwell ;
        RECT 2.930 268.720 343.710 272.240 ;
      LAYER Nwell ;
        RECT 2.930 264.400 343.710 268.720 ;
      LAYER Pwell ;
        RECT 2.930 260.880 343.710 264.400 ;
      LAYER Nwell ;
        RECT 2.930 256.560 343.710 260.880 ;
      LAYER Pwell ;
        RECT 2.930 253.040 343.710 256.560 ;
      LAYER Nwell ;
        RECT 2.930 248.720 343.710 253.040 ;
      LAYER Pwell ;
        RECT 2.930 245.200 343.710 248.720 ;
      LAYER Nwell ;
        RECT 2.930 240.880 343.710 245.200 ;
      LAYER Pwell ;
        RECT 2.930 237.360 343.710 240.880 ;
      LAYER Nwell ;
        RECT 2.930 233.040 343.710 237.360 ;
      LAYER Pwell ;
        RECT 2.930 229.520 343.710 233.040 ;
      LAYER Nwell ;
        RECT 2.930 225.200 343.710 229.520 ;
      LAYER Pwell ;
        RECT 2.930 221.680 343.710 225.200 ;
      LAYER Nwell ;
        RECT 2.930 217.360 343.710 221.680 ;
      LAYER Pwell ;
        RECT 2.930 213.840 343.710 217.360 ;
      LAYER Nwell ;
        RECT 2.930 209.520 343.710 213.840 ;
      LAYER Pwell ;
        RECT 2.930 206.000 343.710 209.520 ;
      LAYER Nwell ;
        RECT 2.930 201.680 343.710 206.000 ;
      LAYER Pwell ;
        RECT 2.930 198.160 343.710 201.680 ;
      LAYER Nwell ;
        RECT 2.930 193.840 343.710 198.160 ;
      LAYER Pwell ;
        RECT 2.930 190.320 343.710 193.840 ;
      LAYER Nwell ;
        RECT 2.930 186.000 343.710 190.320 ;
      LAYER Pwell ;
        RECT 2.930 182.480 343.710 186.000 ;
      LAYER Nwell ;
        RECT 2.930 178.160 343.710 182.480 ;
      LAYER Pwell ;
        RECT 2.930 174.640 343.710 178.160 ;
      LAYER Nwell ;
        RECT 2.930 170.320 343.710 174.640 ;
      LAYER Pwell ;
        RECT 2.930 166.800 343.710 170.320 ;
      LAYER Nwell ;
        RECT 2.930 162.480 343.710 166.800 ;
      LAYER Pwell ;
        RECT 2.930 158.960 343.710 162.480 ;
      LAYER Nwell ;
        RECT 2.930 154.640 343.710 158.960 ;
      LAYER Pwell ;
        RECT 2.930 151.120 343.710 154.640 ;
      LAYER Nwell ;
        RECT 2.930 146.800 343.710 151.120 ;
      LAYER Pwell ;
        RECT 2.930 143.280 343.710 146.800 ;
      LAYER Nwell ;
        RECT 2.930 138.960 343.710 143.280 ;
      LAYER Pwell ;
        RECT 2.930 135.440 343.710 138.960 ;
      LAYER Nwell ;
        RECT 2.930 131.120 343.710 135.440 ;
      LAYER Pwell ;
        RECT 2.930 127.600 343.710 131.120 ;
      LAYER Nwell ;
        RECT 2.930 123.280 343.710 127.600 ;
      LAYER Pwell ;
        RECT 2.930 119.760 343.710 123.280 ;
      LAYER Nwell ;
        RECT 2.930 115.440 343.710 119.760 ;
      LAYER Pwell ;
        RECT 2.930 111.920 343.710 115.440 ;
      LAYER Nwell ;
        RECT 2.930 107.600 343.710 111.920 ;
      LAYER Pwell ;
        RECT 2.930 104.080 343.710 107.600 ;
      LAYER Nwell ;
        RECT 2.930 99.760 343.710 104.080 ;
      LAYER Pwell ;
        RECT 2.930 96.240 343.710 99.760 ;
      LAYER Nwell ;
        RECT 2.930 91.920 343.710 96.240 ;
      LAYER Pwell ;
        RECT 2.930 88.400 343.710 91.920 ;
      LAYER Nwell ;
        RECT 2.930 84.080 343.710 88.400 ;
      LAYER Pwell ;
        RECT 2.930 80.560 343.710 84.080 ;
      LAYER Nwell ;
        RECT 2.930 76.240 343.710 80.560 ;
      LAYER Pwell ;
        RECT 2.930 72.720 343.710 76.240 ;
      LAYER Nwell ;
        RECT 2.930 68.400 343.710 72.720 ;
      LAYER Pwell ;
        RECT 2.930 64.880 343.710 68.400 ;
      LAYER Nwell ;
        RECT 2.930 60.560 343.710 64.880 ;
      LAYER Pwell ;
        RECT 2.930 57.040 343.710 60.560 ;
      LAYER Nwell ;
        RECT 2.930 52.720 343.710 57.040 ;
      LAYER Pwell ;
        RECT 2.930 49.200 343.710 52.720 ;
      LAYER Nwell ;
        RECT 2.930 44.880 343.710 49.200 ;
      LAYER Pwell ;
        RECT 2.930 41.360 343.710 44.880 ;
      LAYER Nwell ;
        RECT 2.930 37.040 343.710 41.360 ;
      LAYER Pwell ;
        RECT 2.930 33.520 343.710 37.040 ;
      LAYER Nwell ;
        RECT 2.930 29.200 343.710 33.520 ;
      LAYER Pwell ;
        RECT 2.930 25.680 343.710 29.200 ;
      LAYER Nwell ;
        RECT 2.930 21.360 343.710 25.680 ;
      LAYER Pwell ;
        RECT 2.930 17.840 343.710 21.360 ;
      LAYER Nwell ;
        RECT 2.930 13.520 343.710 17.840 ;
      LAYER Pwell ;
        RECT 2.930 10.000 343.710 13.520 ;
      LAYER Nwell ;
        RECT 2.930 5.680 343.710 10.000 ;
      LAYER Pwell ;
        RECT 2.930 3.490 343.710 5.680 ;
      LAYER Metal1 ;
        RECT 3.360 3.620 343.280 321.740 ;
      LAYER Metal2 ;
        RECT 5.740 3.730 344.820 322.470 ;
      LAYER Metal3 ;
        RECT 5.690 3.780 344.870 322.420 ;
      LAYER Metal4 ;
        RECT 33.210 324.060 39.590 324.360 ;
        RECT 40.490 324.060 46.870 324.360 ;
        RECT 47.770 324.060 54.150 324.360 ;
        RECT 55.050 324.060 61.430 324.360 ;
        RECT 62.330 324.060 68.710 324.360 ;
        RECT 69.610 324.060 75.990 324.360 ;
        RECT 76.890 324.060 83.270 324.360 ;
        RECT 84.170 324.060 90.550 324.360 ;
        RECT 91.450 324.060 97.830 324.360 ;
        RECT 98.730 324.060 105.110 324.360 ;
        RECT 106.010 324.060 112.390 324.360 ;
        RECT 113.290 324.060 119.670 324.360 ;
        RECT 120.570 324.060 126.950 324.360 ;
        RECT 127.850 324.060 134.230 324.360 ;
        RECT 135.130 324.060 141.510 324.360 ;
        RECT 142.410 324.060 148.790 324.360 ;
        RECT 149.690 324.060 156.070 324.360 ;
        RECT 156.970 324.060 163.350 324.360 ;
        RECT 164.250 324.060 170.630 324.360 ;
        RECT 171.530 324.060 177.910 324.360 ;
        RECT 178.810 324.060 185.190 324.360 ;
        RECT 186.090 324.060 192.470 324.360 ;
        RECT 193.370 324.060 199.750 324.360 ;
        RECT 200.650 324.060 207.030 324.360 ;
        RECT 207.930 324.060 214.310 324.360 ;
        RECT 215.210 324.060 221.590 324.360 ;
        RECT 222.490 324.060 228.870 324.360 ;
        RECT 229.770 324.060 236.150 324.360 ;
        RECT 237.050 324.060 243.430 324.360 ;
        RECT 244.330 324.060 250.710 324.360 ;
        RECT 251.610 324.060 257.990 324.360 ;
        RECT 258.890 324.060 265.270 324.360 ;
        RECT 266.170 324.060 272.550 324.360 ;
        RECT 273.450 324.060 279.830 324.360 ;
        RECT 280.730 324.060 287.110 324.360 ;
        RECT 288.010 324.060 294.390 324.360 ;
        RECT 295.290 324.060 301.670 324.360 ;
        RECT 302.570 324.060 308.950 324.360 ;
        RECT 309.850 324.060 316.230 324.360 ;
        RECT 317.130 324.060 323.510 324.360 ;
        RECT 324.410 324.060 330.790 324.360 ;
        RECT 331.690 324.060 338.070 324.360 ;
        RECT 338.970 324.060 340.900 324.360 ;
        RECT 32.620 322.040 340.900 324.060 ;
        RECT 32.620 6.250 57.450 322.040 ;
        RECT 59.650 6.250 60.750 322.040 ;
        RECT 62.950 6.250 96.320 322.040 ;
        RECT 98.520 6.250 99.620 322.040 ;
        RECT 101.820 6.250 135.190 322.040 ;
        RECT 137.390 6.250 138.490 322.040 ;
        RECT 140.690 6.250 174.060 322.040 ;
        RECT 176.260 6.250 177.360 322.040 ;
        RECT 179.560 6.250 212.930 322.040 ;
        RECT 215.130 6.250 216.230 322.040 ;
        RECT 218.430 6.250 251.800 322.040 ;
        RECT 254.000 6.250 255.100 322.040 ;
        RECT 257.300 6.250 290.670 322.040 ;
        RECT 292.870 6.250 293.970 322.040 ;
        RECT 296.170 6.250 329.540 322.040 ;
        RECT 331.740 6.250 332.840 322.040 ;
        RECT 335.040 6.250 340.900 322.040 ;
  END
END tt_um_a1k0n_nyancat
END LIBRARY

