VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_calonso88_spi_i2c_reg_bank
  CLASS BLOCK ;
  FOREIGN tt_um_calonso88_spi_i2c_reg_bank ;
  ORIGIN 0.000 0.000 ;
  SIZE 346.640 BY 160.720 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 3.620 23.780 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 61.050 3.620 62.650 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.920 3.620 101.520 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.790 3.620 140.390 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 177.660 3.620 179.260 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 216.530 3.620 218.130 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 255.400 3.620 257.000 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 294.270 3.620 295.870 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 333.140 3.620 334.740 157.100 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 3.620 20.480 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 57.750 3.620 59.350 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 96.620 3.620 98.220 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 135.490 3.620 137.090 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 174.360 3.620 175.960 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 213.230 3.620 214.830 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.100 3.620 253.700 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 290.970 3.620 292.570 157.100 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.840 3.620 331.440 157.100 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    PORT
      LAYER Metal4 ;
        RECT 312.890 159.720 313.190 160.720 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 320.170 159.720 320.470 160.720 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 305.610 159.720 305.910 160.720 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 298.330 159.720 298.630 160.720 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 291.050 159.720 291.350 160.720 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 283.770 159.720 284.070 160.720 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 276.490 159.720 276.790 160.720 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 269.210 159.720 269.510 160.720 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 261.930 159.720 262.230 160.720 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 254.650 159.720 254.950 160.720 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 247.370 159.720 247.670 160.720 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 240.090 159.720 240.390 160.720 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 232.810 159.720 233.110 160.720 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 225.530 159.720 225.830 160.720 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 218.250 159.720 218.550 160.720 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    PORT
      LAYER Metal4 ;
        RECT 210.970 159.720 211.270 160.720 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 203.690 159.720 203.990 160.720 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 196.410 159.720 196.710 160.720 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 189.130 159.720 189.430 160.720 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 65.370 159.720 65.670 160.720 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal4 ;
        RECT 58.090 159.720 58.390 160.720 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 50.810 159.720 51.110 160.720 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.099500 ;
    ANTENNADIFFAREA 2.609600 ;
    PORT
      LAYER Metal4 ;
        RECT 43.530 159.720 43.830 160.720 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 36.250 159.720 36.550 160.720 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 28.970 159.720 29.270 160.720 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 21.690 159.720 21.990 160.720 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 14.410 159.720 14.710 160.720 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 123.610 159.720 123.910 160.720 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 116.330 159.720 116.630 160.720 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 109.050 159.720 109.350 160.720 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal4 ;
        RECT 101.770 159.720 102.070 160.720 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 94.490 159.720 94.790 160.720 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 87.210 159.720 87.510 160.720 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 79.930 159.720 80.230 160.720 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 72.650 159.720 72.950 160.720 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 181.850 159.720 182.150 160.720 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 174.570 159.720 174.870 160.720 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 167.290 159.720 167.590 160.720 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 160.010 159.720 160.310 160.720 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 152.730 159.720 153.030 160.720 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 145.450 159.720 145.750 160.720 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 138.170 159.720 138.470 160.720 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal4 ;
        RECT 130.890 159.720 131.190 160.720 ;
    END
  END uo_out[7]
  OBS
      LAYER Nwell ;
        RECT 2.930 154.640 343.710 157.230 ;
      LAYER Pwell ;
        RECT 2.930 151.120 343.710 154.640 ;
      LAYER Nwell ;
        RECT 2.930 146.800 343.710 151.120 ;
      LAYER Pwell ;
        RECT 2.930 143.280 343.710 146.800 ;
      LAYER Nwell ;
        RECT 2.930 138.960 343.710 143.280 ;
      LAYER Pwell ;
        RECT 2.930 135.440 343.710 138.960 ;
      LAYER Nwell ;
        RECT 2.930 131.120 343.710 135.440 ;
      LAYER Pwell ;
        RECT 2.930 127.600 343.710 131.120 ;
      LAYER Nwell ;
        RECT 2.930 123.280 343.710 127.600 ;
      LAYER Pwell ;
        RECT 2.930 119.760 343.710 123.280 ;
      LAYER Nwell ;
        RECT 2.930 115.440 343.710 119.760 ;
      LAYER Pwell ;
        RECT 2.930 111.920 343.710 115.440 ;
      LAYER Nwell ;
        RECT 2.930 107.600 343.710 111.920 ;
      LAYER Pwell ;
        RECT 2.930 104.080 343.710 107.600 ;
      LAYER Nwell ;
        RECT 2.930 99.760 343.710 104.080 ;
      LAYER Pwell ;
        RECT 2.930 96.240 343.710 99.760 ;
      LAYER Nwell ;
        RECT 2.930 91.920 343.710 96.240 ;
      LAYER Pwell ;
        RECT 2.930 88.400 343.710 91.920 ;
      LAYER Nwell ;
        RECT 2.930 84.080 343.710 88.400 ;
      LAYER Pwell ;
        RECT 2.930 80.560 343.710 84.080 ;
      LAYER Nwell ;
        RECT 2.930 76.240 343.710 80.560 ;
      LAYER Pwell ;
        RECT 2.930 72.720 343.710 76.240 ;
      LAYER Nwell ;
        RECT 2.930 68.400 343.710 72.720 ;
      LAYER Pwell ;
        RECT 2.930 64.880 343.710 68.400 ;
      LAYER Nwell ;
        RECT 2.930 60.560 343.710 64.880 ;
      LAYER Pwell ;
        RECT 2.930 57.040 343.710 60.560 ;
      LAYER Nwell ;
        RECT 2.930 52.720 343.710 57.040 ;
      LAYER Pwell ;
        RECT 2.930 49.200 343.710 52.720 ;
      LAYER Nwell ;
        RECT 2.930 44.880 343.710 49.200 ;
      LAYER Pwell ;
        RECT 2.930 41.360 343.710 44.880 ;
      LAYER Nwell ;
        RECT 2.930 37.040 343.710 41.360 ;
      LAYER Pwell ;
        RECT 2.930 33.520 343.710 37.040 ;
      LAYER Nwell ;
        RECT 2.930 29.200 343.710 33.520 ;
      LAYER Pwell ;
        RECT 2.930 25.680 343.710 29.200 ;
      LAYER Nwell ;
        RECT 2.930 21.360 343.710 25.680 ;
      LAYER Pwell ;
        RECT 2.930 17.840 343.710 21.360 ;
      LAYER Nwell ;
        RECT 2.930 13.520 343.710 17.840 ;
      LAYER Pwell ;
        RECT 2.930 10.000 343.710 13.520 ;
      LAYER Nwell ;
        RECT 2.930 5.680 343.710 10.000 ;
      LAYER Pwell ;
        RECT 2.930 3.490 343.710 5.680 ;
      LAYER Metal1 ;
        RECT 3.360 3.620 343.280 157.100 ;
      LAYER Metal2 ;
        RECT 15.260 3.730 340.900 158.390 ;
      LAYER Metal3 ;
        RECT 14.370 3.780 339.830 158.340 ;
      LAYER Metal4 ;
        RECT 15.010 159.420 21.390 159.720 ;
        RECT 22.290 159.420 28.670 159.720 ;
        RECT 29.570 159.420 35.950 159.720 ;
        RECT 36.850 159.420 43.230 159.720 ;
        RECT 44.130 159.420 50.510 159.720 ;
        RECT 51.410 159.420 57.790 159.720 ;
        RECT 58.690 159.420 65.070 159.720 ;
        RECT 65.970 159.420 72.350 159.720 ;
        RECT 73.250 159.420 79.630 159.720 ;
        RECT 80.530 159.420 86.910 159.720 ;
        RECT 87.810 159.420 94.190 159.720 ;
        RECT 95.090 159.420 101.470 159.720 ;
        RECT 102.370 159.420 108.750 159.720 ;
        RECT 109.650 159.420 116.030 159.720 ;
        RECT 116.930 159.420 123.310 159.720 ;
        RECT 124.210 159.420 130.590 159.720 ;
        RECT 131.490 159.420 137.870 159.720 ;
        RECT 138.770 159.420 145.150 159.720 ;
        RECT 146.050 159.420 152.430 159.720 ;
        RECT 153.330 159.420 159.710 159.720 ;
        RECT 160.610 159.420 166.990 159.720 ;
        RECT 167.890 159.420 174.270 159.720 ;
        RECT 175.170 159.420 181.550 159.720 ;
        RECT 182.450 159.420 188.830 159.720 ;
        RECT 189.730 159.420 196.110 159.720 ;
        RECT 197.010 159.420 203.390 159.720 ;
        RECT 204.290 159.420 210.670 159.720 ;
        RECT 211.570 159.420 217.950 159.720 ;
        RECT 218.850 159.420 225.230 159.720 ;
        RECT 226.130 159.420 232.510 159.720 ;
        RECT 233.410 159.420 239.790 159.720 ;
        RECT 240.690 159.420 247.070 159.720 ;
        RECT 247.970 159.420 254.350 159.720 ;
        RECT 255.250 159.420 261.630 159.720 ;
        RECT 262.530 159.420 268.910 159.720 ;
        RECT 269.810 159.420 276.190 159.720 ;
        RECT 277.090 159.420 283.470 159.720 ;
        RECT 284.370 159.420 290.750 159.720 ;
        RECT 291.650 159.420 298.030 159.720 ;
        RECT 298.930 159.420 305.310 159.720 ;
        RECT 306.210 159.420 312.590 159.720 ;
        RECT 313.490 159.420 319.870 159.720 ;
        RECT 14.420 157.400 320.460 159.420 ;
        RECT 14.420 33.690 18.580 157.400 ;
        RECT 20.780 33.690 21.880 157.400 ;
        RECT 24.080 33.690 57.450 157.400 ;
        RECT 59.650 33.690 60.750 157.400 ;
        RECT 62.950 33.690 96.320 157.400 ;
        RECT 98.520 33.690 99.620 157.400 ;
        RECT 101.820 33.690 135.190 157.400 ;
        RECT 137.390 33.690 138.490 157.400 ;
        RECT 140.690 33.690 174.060 157.400 ;
        RECT 176.260 33.690 177.360 157.400 ;
        RECT 179.560 33.690 212.930 157.400 ;
        RECT 215.130 33.690 216.230 157.400 ;
        RECT 218.430 33.690 251.800 157.400 ;
        RECT 254.000 33.690 255.100 157.400 ;
        RECT 257.300 33.690 290.670 157.400 ;
        RECT 292.870 33.690 293.970 157.400 ;
        RECT 296.170 33.690 320.460 157.400 ;
  END
END tt_um_calonso88_spi_i2c_reg_bank
END LIBRARY

