VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_rejunity_vga_test01
  CLASS BLOCK ;
  FOREIGN tt_um_rejunity_vga_test01 ;
  ORIGIN 0.000 0.000 ;
  SIZE 711.200 BY 325.360 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 22.180 4.740 23.780 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 61.050 4.740 62.650 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.920 4.740 101.520 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 138.790 4.740 140.390 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 177.660 4.740 179.260 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 216.530 4.740 218.130 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 255.400 4.740 257.000 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 294.270 4.740 295.870 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 333.140 4.740 334.740 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 372.010 4.740 373.610 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 410.880 4.740 412.480 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 449.750 4.740 451.350 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 488.620 4.740 490.220 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 527.490 4.740 529.090 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 566.360 4.740 567.960 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.230 4.740 606.830 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 644.100 4.740 645.700 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 682.970 4.740 684.570 317.820 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.880 4.740 20.480 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 57.750 4.740 59.350 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 96.620 4.740 98.220 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 135.490 4.740 137.090 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 174.360 4.740 175.960 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 213.230 4.740 214.830 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.100 4.740 253.700 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 290.970 4.740 292.570 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.840 4.740 331.440 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 368.710 4.740 370.310 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 407.580 4.740 409.180 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 446.450 4.740 448.050 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 485.320 4.740 486.920 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 524.190 4.740 525.790 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 563.060 4.740 564.660 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 601.930 4.740 603.530 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 640.800 4.740 642.400 317.820 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 679.670 4.740 681.270 317.820 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.823999 ;
    PORT
      LAYER Metal4 ;
        RECT 331.090 324.360 331.390 325.360 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 338.370 324.360 338.670 325.360 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 323.810 324.360 324.110 325.360 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 316.530 324.360 316.830 325.360 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 309.250 324.360 309.550 325.360 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 301.970 324.360 302.270 325.360 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 294.690 324.360 294.990 325.360 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 287.410 324.360 287.710 325.360 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 280.130 324.360 280.430 325.360 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 272.850 324.360 273.150 325.360 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 265.570 324.360 265.870 325.360 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 258.290 324.360 258.590 325.360 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 251.010 324.360 251.310 325.360 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 243.730 324.360 244.030 325.360 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 236.450 324.360 236.750 325.360 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 229.170 324.360 229.470 325.360 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 221.890 324.360 222.190 325.360 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 214.610 324.360 214.910 325.360 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 207.330 324.360 207.630 325.360 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 83.570 324.360 83.870 325.360 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 76.290 324.360 76.590 325.360 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 69.010 324.360 69.310 325.360 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 61.730 324.360 62.030 325.360 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 54.450 324.360 54.750 325.360 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 47.170 324.360 47.470 325.360 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 39.890 324.360 40.190 325.360 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.396000 ;
    PORT
      LAYER Metal4 ;
        RECT 32.610 324.360 32.910 325.360 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal4 ;
        RECT 141.810 324.360 142.110 325.360 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal4 ;
        RECT 134.530 324.360 134.830 325.360 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal4 ;
        RECT 127.250 324.360 127.550 325.360 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal4 ;
        RECT 119.970 324.360 120.270 325.360 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal4 ;
        RECT 112.690 324.360 112.990 325.360 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal4 ;
        RECT 105.410 324.360 105.710 325.360 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.821000 ;
    PORT
      LAYER Metal4 ;
        RECT 98.130 324.360 98.430 325.360 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 11.948999 ;
    ANTENNADIFFAREA 3.276000 ;
    PORT
      LAYER Metal4 ;
        RECT 90.850 324.360 91.150 325.360 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal4 ;
        RECT 200.050 324.360 200.350 325.360 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal4 ;
        RECT 192.770 324.360 193.070 325.360 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal4 ;
        RECT 185.490 324.360 185.790 325.360 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal4 ;
        RECT 178.210 324.360 178.510 325.360 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal4 ;
        RECT 170.930 324.360 171.230 325.360 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal4 ;
        RECT 163.650 324.360 163.950 325.360 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal4 ;
        RECT 156.370 324.360 156.670 325.360 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.638000 ;
    PORT
      LAYER Metal4 ;
        RECT 149.090 324.360 149.390 325.360 ;
    END
  END uo_out[7]
  OBS
      LAYER Pwell ;
        RECT 0.430 315.255 710.770 317.950 ;
      LAYER Nwell ;
        RECT 0.430 309.705 710.770 315.255 ;
      LAYER Pwell ;
        RECT 0.430 305.175 710.770 309.705 ;
      LAYER Nwell ;
        RECT 0.430 299.625 710.770 305.175 ;
      LAYER Pwell ;
        RECT 0.430 295.095 710.770 299.625 ;
      LAYER Nwell ;
        RECT 0.430 289.545 710.770 295.095 ;
      LAYER Pwell ;
        RECT 0.430 285.015 710.770 289.545 ;
      LAYER Nwell ;
        RECT 0.430 279.465 710.770 285.015 ;
      LAYER Pwell ;
        RECT 0.430 274.935 710.770 279.465 ;
      LAYER Nwell ;
        RECT 0.430 269.385 710.770 274.935 ;
      LAYER Pwell ;
        RECT 0.430 264.855 710.770 269.385 ;
      LAYER Nwell ;
        RECT 0.430 259.305 710.770 264.855 ;
      LAYER Pwell ;
        RECT 0.430 254.775 710.770 259.305 ;
      LAYER Nwell ;
        RECT 0.430 249.225 710.770 254.775 ;
      LAYER Pwell ;
        RECT 0.430 244.695 710.770 249.225 ;
      LAYER Nwell ;
        RECT 0.430 239.145 710.770 244.695 ;
      LAYER Pwell ;
        RECT 0.430 234.615 710.770 239.145 ;
      LAYER Nwell ;
        RECT 0.430 229.065 710.770 234.615 ;
      LAYER Pwell ;
        RECT 0.430 224.535 710.770 229.065 ;
      LAYER Nwell ;
        RECT 0.430 218.985 710.770 224.535 ;
      LAYER Pwell ;
        RECT 0.430 214.455 710.770 218.985 ;
      LAYER Nwell ;
        RECT 0.430 208.905 710.770 214.455 ;
      LAYER Pwell ;
        RECT 0.430 204.375 710.770 208.905 ;
      LAYER Nwell ;
        RECT 0.430 198.825 710.770 204.375 ;
      LAYER Pwell ;
        RECT 0.430 194.295 710.770 198.825 ;
      LAYER Nwell ;
        RECT 0.430 188.745 710.770 194.295 ;
      LAYER Pwell ;
        RECT 0.430 184.215 710.770 188.745 ;
      LAYER Nwell ;
        RECT 0.430 178.665 710.770 184.215 ;
      LAYER Pwell ;
        RECT 0.430 174.135 710.770 178.665 ;
      LAYER Nwell ;
        RECT 0.430 168.585 710.770 174.135 ;
      LAYER Pwell ;
        RECT 0.430 164.055 710.770 168.585 ;
      LAYER Nwell ;
        RECT 0.430 158.505 710.770 164.055 ;
      LAYER Pwell ;
        RECT 0.430 153.975 710.770 158.505 ;
      LAYER Nwell ;
        RECT 0.430 148.425 710.770 153.975 ;
      LAYER Pwell ;
        RECT 0.430 143.895 710.770 148.425 ;
      LAYER Nwell ;
        RECT 0.430 138.345 710.770 143.895 ;
      LAYER Pwell ;
        RECT 0.430 133.815 710.770 138.345 ;
      LAYER Nwell ;
        RECT 0.430 128.265 710.770 133.815 ;
      LAYER Pwell ;
        RECT 0.430 123.735 710.770 128.265 ;
      LAYER Nwell ;
        RECT 0.430 118.185 710.770 123.735 ;
      LAYER Pwell ;
        RECT 0.430 113.655 710.770 118.185 ;
      LAYER Nwell ;
        RECT 0.430 108.105 710.770 113.655 ;
      LAYER Pwell ;
        RECT 0.430 103.575 710.770 108.105 ;
      LAYER Nwell ;
        RECT 0.430 98.025 710.770 103.575 ;
      LAYER Pwell ;
        RECT 0.430 93.495 710.770 98.025 ;
      LAYER Nwell ;
        RECT 0.430 87.945 710.770 93.495 ;
      LAYER Pwell ;
        RECT 0.430 83.415 710.770 87.945 ;
      LAYER Nwell ;
        RECT 0.430 77.865 710.770 83.415 ;
      LAYER Pwell ;
        RECT 0.430 73.335 710.770 77.865 ;
      LAYER Nwell ;
        RECT 0.430 67.785 710.770 73.335 ;
      LAYER Pwell ;
        RECT 0.430 63.255 710.770 67.785 ;
      LAYER Nwell ;
        RECT 0.430 57.705 710.770 63.255 ;
      LAYER Pwell ;
        RECT 0.430 53.175 710.770 57.705 ;
      LAYER Nwell ;
        RECT 0.430 47.625 710.770 53.175 ;
      LAYER Pwell ;
        RECT 0.430 43.095 710.770 47.625 ;
      LAYER Nwell ;
        RECT 0.430 37.545 710.770 43.095 ;
      LAYER Pwell ;
        RECT 0.430 33.015 710.770 37.545 ;
      LAYER Nwell ;
        RECT 0.430 27.465 710.770 33.015 ;
      LAYER Pwell ;
        RECT 0.430 22.935 710.770 27.465 ;
      LAYER Nwell ;
        RECT 0.430 17.385 710.770 22.935 ;
      LAYER Pwell ;
        RECT 0.430 12.855 710.770 17.385 ;
      LAYER Nwell ;
        RECT 0.430 7.305 710.770 12.855 ;
      LAYER Pwell ;
        RECT 0.430 4.610 710.770 7.305 ;
      LAYER Metal1 ;
        RECT 3.360 4.590 707.840 317.970 ;
      LAYER Metal2 ;
        RECT 5.180 4.850 684.430 320.230 ;
      LAYER Metal3 ;
        RECT 5.130 4.900 684.480 320.180 ;
      LAYER Metal4 ;
        RECT 33.210 324.060 39.590 324.360 ;
        RECT 40.490 324.060 46.870 324.360 ;
        RECT 47.770 324.060 54.150 324.360 ;
        RECT 55.050 324.060 61.430 324.360 ;
        RECT 62.330 324.060 68.710 324.360 ;
        RECT 69.610 324.060 75.990 324.360 ;
        RECT 76.890 324.060 83.270 324.360 ;
        RECT 84.170 324.060 90.550 324.360 ;
        RECT 91.450 324.060 97.830 324.360 ;
        RECT 98.730 324.060 105.110 324.360 ;
        RECT 106.010 324.060 112.390 324.360 ;
        RECT 113.290 324.060 119.670 324.360 ;
        RECT 120.570 324.060 126.950 324.360 ;
        RECT 127.850 324.060 134.230 324.360 ;
        RECT 135.130 324.060 141.510 324.360 ;
        RECT 142.410 324.060 148.790 324.360 ;
        RECT 149.690 324.060 156.070 324.360 ;
        RECT 156.970 324.060 163.350 324.360 ;
        RECT 164.250 324.060 170.630 324.360 ;
        RECT 171.530 324.060 177.910 324.360 ;
        RECT 178.810 324.060 185.190 324.360 ;
        RECT 186.090 324.060 192.470 324.360 ;
        RECT 193.370 324.060 199.750 324.360 ;
        RECT 200.650 324.060 207.030 324.360 ;
        RECT 207.930 324.060 214.310 324.360 ;
        RECT 215.210 324.060 221.590 324.360 ;
        RECT 222.490 324.060 228.870 324.360 ;
        RECT 229.770 324.060 236.150 324.360 ;
        RECT 237.050 324.060 243.430 324.360 ;
        RECT 244.330 324.060 250.710 324.360 ;
        RECT 251.610 324.060 257.990 324.360 ;
        RECT 258.890 324.060 265.270 324.360 ;
        RECT 266.170 324.060 272.550 324.360 ;
        RECT 273.450 324.060 279.830 324.360 ;
        RECT 280.730 324.060 287.110 324.360 ;
        RECT 288.010 324.060 294.390 324.360 ;
        RECT 295.290 324.060 301.670 324.360 ;
        RECT 302.570 324.060 308.950 324.360 ;
        RECT 309.850 324.060 316.230 324.360 ;
        RECT 317.130 324.060 323.510 324.360 ;
        RECT 324.410 324.060 330.790 324.360 ;
        RECT 331.690 324.060 338.070 324.360 ;
        RECT 338.970 324.060 590.660 324.360 ;
        RECT 32.620 318.120 590.660 324.060 ;
        RECT 32.620 21.930 57.450 318.120 ;
        RECT 59.650 21.930 60.750 318.120 ;
        RECT 62.950 21.930 96.320 318.120 ;
        RECT 98.520 21.930 99.620 318.120 ;
        RECT 101.820 21.930 135.190 318.120 ;
        RECT 137.390 21.930 138.490 318.120 ;
        RECT 140.690 21.930 174.060 318.120 ;
        RECT 176.260 21.930 177.360 318.120 ;
        RECT 179.560 21.930 212.930 318.120 ;
        RECT 215.130 21.930 216.230 318.120 ;
        RECT 218.430 21.930 251.800 318.120 ;
        RECT 254.000 21.930 255.100 318.120 ;
        RECT 257.300 21.930 290.670 318.120 ;
        RECT 292.870 21.930 293.970 318.120 ;
        RECT 296.170 21.930 329.540 318.120 ;
        RECT 331.740 21.930 332.840 318.120 ;
        RECT 335.040 21.930 368.410 318.120 ;
        RECT 370.610 21.930 371.710 318.120 ;
        RECT 373.910 21.930 407.280 318.120 ;
        RECT 409.480 21.930 410.580 318.120 ;
        RECT 412.780 21.930 446.150 318.120 ;
        RECT 448.350 21.930 449.450 318.120 ;
        RECT 451.650 21.930 485.020 318.120 ;
        RECT 487.220 21.930 488.320 318.120 ;
        RECT 490.520 21.930 523.890 318.120 ;
        RECT 526.090 21.930 527.190 318.120 ;
        RECT 529.390 21.930 562.760 318.120 ;
        RECT 564.960 21.930 566.060 318.120 ;
        RECT 568.260 21.930 590.660 318.120 ;
  END
END tt_um_rejunity_vga_test01
END LIBRARY

