module tt_um_rejunity_vga_test01 (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire \center_x[0] ;
 wire \center_x[1] ;
 wire \center_x[2] ;
 wire \center_x[3] ;
 wire \center_x[4] ;
 wire \center_x[5] ;
 wire \center_y[0] ;
 wire \dot2[0] ;
 wire \dot2[1] ;
 wire \dot2[2] ;
 wire \dot2[3] ;
 wire \dot2[4] ;
 wire \dot2[5] ;
 wire \dot2[6] ;
 wire \dot2[7] ;
 wire \dot[0] ;
 wire \dot[1] ;
 wire \dot[2] ;
 wire \dot[3] ;
 wire \dot[4] ;
 wire \dot[5] ;
 wire \dot[6] ;
 wire \dot[7] ;
 wire \dot__t[0] ;
 wire \dot__t[1] ;
 wire \dot__t[2] ;
 wire \dot__t[3] ;
 wire \dot__t[4] ;
 wire \dot__t[5] ;
 wire \dot__t[6] ;
 wire \dot__t[7] ;
 wire \frame_counter[7] ;
 wire \frame_counter[8] ;
 wire \frame_counter[9] ;
 wire frame_counter_frac;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire noise;
 wire \noise_counter[0] ;
 wire \noise_counter[1] ;
 wire \noise_counter[2] ;
 wire note;
 wire note2;
 wire \note2_counter[0] ;
 wire \note2_counter[1] ;
 wire \note2_counter[2] ;
 wire \note2_counter[3] ;
 wire \note2_counter[4] ;
 wire \note2_counter[5] ;
 wire \note2_counter[6] ;
 wire \note2_counter[7] ;
 wire \note2_counter[8] ;
 wire \note2_freq[0] ;
 wire \note2_freq[1] ;
 wire \note2_freq[3] ;
 wire \note2_freq[4] ;
 wire \note2_freq[5] ;
 wire \note2_freq[6] ;
 wire \note2_freq[7] ;
 wire \note2_freq[8] ;
 wire \note_counter[0] ;
 wire \note_counter[1] ;
 wire \note_counter[2] ;
 wire \note_counter[3] ;
 wire \note_counter[4] ;
 wire \note_counter[5] ;
 wire \note_counter[6] ;
 wire \note_counter[7] ;
 wire \note_freq[0] ;
 wire \note_freq[1] ;
 wire \note_freq[2] ;
 wire \note_freq[4] ;
 wire \note_freq[5] ;
 wire \note_freq[6] ;
 wire \note_freq[7] ;
 wire \p_p[0] ;
 wire \p_p[1] ;
 wire \p_p[2] ;
 wire \p_p[3] ;
 wire \p_p[4] ;
 wire \p_p[5] ;
 wire \p_p[6] ;
 wire \p_p[7] ;
 wire \p_p__t[0] ;
 wire \p_p__t[1] ;
 wire \p_p__t[2] ;
 wire \p_p__t[3] ;
 wire \p_p__t[4] ;
 wire \p_p__t[5] ;
 wire \p_p__t[6] ;
 wire \p_p__t[7] ;
 wire \pp_x_sq[0] ;
 wire \pp_x_sq[10] ;
 wire \pp_x_sq[11] ;
 wire \pp_x_sq[12] ;
 wire \pp_x_sq[13] ;
 wire \pp_x_sq[14] ;
 wire \pp_x_sq[15] ;
 wire \pp_x_sq[2] ;
 wire \pp_x_sq[3] ;
 wire \pp_x_sq[4] ;
 wire \pp_x_sq[5] ;
 wire \pp_x_sq[6] ;
 wire \pp_x_sq[7] ;
 wire \pp_x_sq[8] ;
 wire \pp_x_sq[9] ;
 wire \pp_x_sq__t[10] ;
 wire \pp_x_sq__t[11] ;
 wire \pp_x_sq__t[12] ;
 wire \pp_x_sq__t[13] ;
 wire \pp_x_sq__t[14] ;
 wire \pp_x_sq__t[15] ;
 wire \pp_x_sq__t[2] ;
 wire \pp_x_sq__t[3] ;
 wire \pp_x_sq__t[4] ;
 wire \pp_x_sq__t[5] ;
 wire \pp_x_sq__t[6] ;
 wire \pp_x_sq__t[7] ;
 wire \pp_x_sq__t[8] ;
 wire \pp_x_sq__t[9] ;
 wire \ppp_x[0] ;
 wire \ppp_x[1] ;
 wire \ppp_x[2] ;
 wire \ppp_x[3] ;
 wire \ppp_x[4] ;
 wire \ppp_x[5] ;
 wire \ppp_x[6] ;
 wire \ppp_x[7] ;
 wire \ppp_y[0] ;
 wire \ppp_y[1] ;
 wire \ppp_y[2] ;
 wire \ppp_y[3] ;
 wire \ppp_y[4] ;
 wire \ppp_y[5] ;
 wire \ppp_y[6] ;
 wire \ppp_y[7] ;
 wire \ppp_y__t[0] ;
 wire \ppp_y__t[1] ;
 wire \ppp_y__t[2] ;
 wire \ppp_y__t[3] ;
 wire \ppp_y__t[4] ;
 wire \ppp_y__t[5] ;
 wire \ppp_y__t[6] ;
 wire \ppp_y__t[7] ;
 wire \r1[0] ;
 wire \r1[10] ;
 wire \r1[11] ;
 wire \r1[12] ;
 wire \r1[13] ;
 wire \r1[14] ;
 wire \r1[15] ;
 wire \r1[16] ;
 wire \r1[17] ;
 wire \r1[1] ;
 wire \r1[2] ;
 wire \r1[3] ;
 wire \r1[4] ;
 wire \r1[5] ;
 wire \r1[6] ;
 wire \r1[7] ;
 wire \r1[8] ;
 wire \r1[9] ;
 wire \r2[0] ;
 wire \r2[10] ;
 wire \r2[11] ;
 wire \r2[12] ;
 wire \r2[13] ;
 wire \r2[14] ;
 wire \r2[15] ;
 wire \r2[16] ;
 wire \r2[17] ;
 wire \r2[18] ;
 wire \r2[1] ;
 wire \r2[2] ;
 wire \r2[3] ;
 wire \r2[4] ;
 wire \r2[5] ;
 wire \r2[6] ;
 wire \r2[7] ;
 wire \r2[8] ;
 wire \r2[9] ;
 wire \r[0] ;
 wire \r[10] ;
 wire \r[11] ;
 wire \r[12] ;
 wire \r[13] ;
 wire \r[14] ;
 wire \r[15] ;
 wire \r[16] ;
 wire \r[17] ;
 wire \r[18] ;
 wire \r[19] ;
 wire \r[1] ;
 wire \r[2] ;
 wire \r[3] ;
 wire \r[4] ;
 wire \r[5] ;
 wire \r[6] ;
 wire \r[7] ;
 wire \r[8] ;
 wire \r[9] ;
 wire \r__t[0] ;
 wire \r__t[10] ;
 wire \r__t[11] ;
 wire \r__t[12] ;
 wire \r__t[13] ;
 wire \r__t[14] ;
 wire \r__t[15] ;
 wire \r__t[16] ;
 wire \r__t[17] ;
 wire \r__t[18] ;
 wire \r__t[19] ;
 wire \r__t[1] ;
 wire \r__t[2] ;
 wire \r__t[3] ;
 wire \r__t[4] ;
 wire \r__t[5] ;
 wire \r__t[6] ;
 wire \r__t[7] ;
 wire \r__t[8] ;
 wire \r__t[9] ;
 wire \title_r[0] ;
 wire \title_r[10] ;
 wire \title_r[11] ;
 wire \title_r[12] ;
 wire \title_r[13] ;
 wire \title_r[1] ;
 wire \title_r[2] ;
 wire \title_r[3] ;
 wire \title_r[4] ;
 wire \title_r[5] ;
 wire \title_r[6] ;
 wire \title_r[7] ;
 wire \title_r[8] ;
 wire \title_r[9] ;
 wire \title_r_pixels_in_scanline[0] ;
 wire \title_r_pixels_in_scanline[1] ;
 wire \title_r_pixels_in_scanline[2] ;
 wire \title_r_pixels_in_scanline[3] ;
 wire \title_r_pixels_in_scanline[4] ;
 wire \title_r_pixels_in_scanline[5] ;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire clknet_leaf_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 gf180mcu_fd_sc_mcu9t5v0__inv_1 _3082_ (.I(\title_r[11] ),
    .ZN(_2534_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3083_ (.I(\title_r[10] ),
    .ZN(_2535_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3084_ (.I(\title_r[9] ),
    .ZN(_2536_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _3085_ (.I(\title_r[8] ),
    .ZN(_2537_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3086_ (.I(\title_r[7] ),
    .ZN(_2538_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3087_ (.I(\title_r[6] ),
    .ZN(_2539_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3088_ (.I(\title_r[4] ),
    .ZN(_2540_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3089_ (.I(\title_r[3] ),
    .ZN(_2541_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3090_ (.I(\title_r[2] ),
    .ZN(_2542_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _3091_ (.I(net111),
    .ZN(_2543_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3092_ (.I(\frame_counter[8] ),
    .ZN(_2544_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _3093_ (.I(\frame_counter[7] ),
    .ZN(_2545_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3094_ (.I(net115),
    .ZN(_2546_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3095_ (.I(net120),
    .ZN(_2547_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _3096_ (.I(net125),
    .ZN(_2548_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _3097_ (.I(net129),
    .ZN(_2549_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _3098_ (.I(net131),
    .ZN(_2550_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _3099_ (.I(net136),
    .ZN(_2551_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _3100_ (.I(net148),
    .ZN(_2552_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3101_ (.I(note),
    .ZN(_2553_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3102_ (.I(\note_counter[7] ),
    .ZN(_2554_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3103_ (.I(\note_counter[2] ),
    .ZN(_2555_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3104_ (.I(\note_counter[0] ),
    .ZN(_2556_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3105_ (.I(\note2_counter[8] ),
    .ZN(_2557_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3106_ (.I(\note2_counter[7] ),
    .ZN(_2558_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3107_ (.I(\note2_counter[6] ),
    .ZN(_2559_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3108_ (.I(\note2_counter[5] ),
    .ZN(_2560_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3109_ (.I(\note2_counter[4] ),
    .ZN(_2561_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3110_ (.I(\note2_counter[3] ),
    .ZN(_2562_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3111_ (.I(\note2_counter[1] ),
    .ZN(_2563_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3112_ (.I(\note2_counter[0] ),
    .ZN(_2564_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3113_ (.I(\title_r[13] ),
    .ZN(_2565_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _3114_ (.I(\hvsync_gen.vpos[0] ),
    .ZN(_2566_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3115_ (.I(\hvsync_gen.hpos[1] ),
    .ZN(_2567_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3116_ (.I(\hvsync_gen.hpos[0] ),
    .ZN(_2568_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3117_ (.I(net161),
    .ZN(_2569_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3118_ (.I(net162),
    .ZN(_2570_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _3119_ (.I(net158),
    .ZN(_2571_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _3120_ (.I(net155),
    .ZN(_2572_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _3121_ (.I(\hvsync_gen.hpos[7] ),
    .ZN(_2573_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _3122_ (.I(net152),
    .ZN(_2574_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _3123_ (.I(\hvsync_gen.hpos[9] ),
    .ZN(_2575_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _3124_ (.I(\hvsync_gen.hpos[8] ),
    .ZN(_2576_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _3125_ (.I(\hvsync_gen.vpos[1] ),
    .ZN(_2577_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3126_ (.I(net97),
    .ZN(_2578_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3127_ (.I(net94),
    .ZN(_2579_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _3128_ (.I(net91),
    .ZN(_2580_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3129_ (.I(\hvsync_gen.vpos[7] ),
    .ZN(_2581_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3130_ (.I(\hvsync_gen.vpos[8] ),
    .ZN(_2582_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _3131_ (.I(\hvsync_gen.vpos[9] ),
    .ZN(_2583_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3132_ (.I(net169),
    .ZN(_2584_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3133_ (.I(\note2_freq[8] ),
    .ZN(_2585_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3134_ (.I(\note_freq[6] ),
    .ZN(_2586_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3135_ (.I(\note_freq[5] ),
    .ZN(_2587_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3136_ (.I(\note_freq[4] ),
    .ZN(_2588_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3137_ (.I(\note_freq[1] ),
    .ZN(_2589_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3138_ (.I(net107),
    .ZN(_2590_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3139_ (.I(\title_r_pixels_in_scanline[2] ),
    .ZN(_2591_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3140_ (.I(\title_r_pixels_in_scanline[0] ),
    .ZN(_2592_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3141_ (.I(net103),
    .ZN(_2593_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3142_ (.I(\ppp_y[6] ),
    .ZN(_2594_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3143_ (.I(net99),
    .ZN(_2595_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3144_ (.I(net89),
    .ZN(_2596_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _3145_ (.I(\r2[1] ),
    .ZN(_2597_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3146_ (.I(\r2[2] ),
    .ZN(_2598_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3147_ (.I(\r2[3] ),
    .ZN(_2599_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3148_ (.I(\r2[4] ),
    .ZN(_2600_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3149_ (.I(\r2[5] ),
    .ZN(_2601_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3150_ (.I(\r2[7] ),
    .ZN(_2602_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3151_ (.I(\r2[8] ),
    .ZN(_2603_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3152_ (.I(\r2[10] ),
    .ZN(_2604_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3153_ (.I(\r2[12] ),
    .ZN(_2605_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _3154_ (.I(\r2[13] ),
    .ZN(_2606_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3155_ (.I(\r2[14] ),
    .ZN(_2607_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3156_ (.I(\r2[17] ),
    .ZN(_2608_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _3157_ (.I(\r1[0] ),
    .ZN(_2609_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _3158_ (.I(\r1[1] ),
    .ZN(_2610_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3159_ (.I(\r1[2] ),
    .ZN(_2611_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3160_ (.I(\r1[3] ),
    .ZN(_2612_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _3161_ (.I(\r1[4] ),
    .ZN(_2613_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3162_ (.I(\r1[6] ),
    .ZN(_2614_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _3163_ (.I(\r1[7] ),
    .ZN(_2615_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3164_ (.I(\r1[8] ),
    .ZN(_2616_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3165_ (.I(\r1[12] ),
    .ZN(_2617_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3166_ (.I(\r1[16] ),
    .ZN(_2618_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3167_ (.I(net106),
    .ZN(_2619_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3168_ (.I(net105),
    .ZN(_2620_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3169_ (.I(\dot[4] ),
    .ZN(_2621_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3170_ (.A1(_2579_),
    .A2(net92),
    .ZN(_2622_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3171_ (.A1(\hvsync_gen.vpos[8] ),
    .A2(_2583_),
    .ZN(_2623_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _3172_ (.A1(\hvsync_gen.vpos[1] ),
    .A2(net95),
    .A3(_2578_),
    .A4(net93),
    .ZN(_2624_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_1 _3173_ (.A1(_2581_),
    .A2(_2622_),
    .A3(_2623_),
    .A4(_2624_),
    .ZN(_0011_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3174_ (.A1(_2573_),
    .A2(\hvsync_gen.hpos[8] ),
    .ZN(_2625_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3175_ (.A1(_2573_),
    .A2(_2575_),
    .A3(\hvsync_gen.hpos[8] ),
    .ZN(_2626_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3176_ (.A1(\hvsync_gen.hpos[9] ),
    .A2(_2625_),
    .ZN(_2627_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_1 _3177_ (.A1(_2571_),
    .A2(_2572_),
    .A3(_2573_),
    .A4(_2574_),
    .ZN(_2628_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3178_ (.A1(net155),
    .A2(net153),
    .ZN(_2629_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _3179_ (.A1(_2571_),
    .A2(_2629_),
    .B(_2628_),
    .C(_2627_),
    .ZN(_0010_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3180_ (.A1(net137),
    .A2(\hvsync_gen.hpos[0] ),
    .ZN(_2630_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3181_ (.A1(net142),
    .A2(\hvsync_gen.hpos[0] ),
    .Z(_2631_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3182_ (.A1(\hvsync_gen.vpos[0] ),
    .A2(net81),
    .ZN(_2632_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3183_ (.A1(net111),
    .A2(_2545_),
    .ZN(_2633_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _3184_ (.A1(net111),
    .A2(\frame_counter[8] ),
    .A3(_2545_),
    .ZN(_2634_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3185_ (.A1(_2543_),
    .A2(_2544_),
    .A3(\frame_counter[7] ),
    .ZN(_2635_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3186_ (.A1(net111),
    .A2(_2545_),
    .ZN(_2636_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _3187_ (.A1(_2543_),
    .A2(_2544_),
    .A3(\frame_counter[7] ),
    .ZN(_2637_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3188_ (.A1(net111),
    .A2(\frame_counter[8] ),
    .A3(_2545_),
    .ZN(_2638_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3189_ (.A1(_2634_),
    .A2(_2637_),
    .ZN(_2639_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _3190_ (.A1(\r[11] ),
    .A2(_2632_),
    .Z(_2640_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3191_ (.A1(\r[11] ),
    .A2(_2632_),
    .B(net60),
    .ZN(_2641_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3192_ (.A1(\ppp_x[0] ),
    .A2(\p_p[0] ),
    .ZN(_2642_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _3193_ (.A1(_2640_),
    .A2(_2641_),
    .B1(_2642_),
    .B2(net60),
    .ZN(\ppp_y__t[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3194_ (.A1(\ppp_x[1] ),
    .A2(\p_p[1] ),
    .ZN(_2643_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3195_ (.A1(\ppp_x[1] ),
    .A2(\p_p[1] ),
    .Z(_2644_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3196_ (.A1(\ppp_x[0] ),
    .A2(\p_p[0] ),
    .B(_2644_),
    .ZN(_2645_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3197_ (.A1(\ppp_x[0] ),
    .A2(\p_p[0] ),
    .A3(_2644_),
    .ZN(_2646_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3198_ (.A1(net60),
    .A2(_2646_),
    .ZN(_2647_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3199_ (.A1(net130),
    .A2(_2567_),
    .ZN(_2648_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3200_ (.A1(net130),
    .A2(\hvsync_gen.hpos[1] ),
    .Z(_2649_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3201_ (.A1(net137),
    .A2(_2568_),
    .B(_2649_),
    .ZN(_2650_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _3202_ (.A1(net137),
    .A2(_2568_),
    .A3(_2649_),
    .Z(_2651_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3203_ (.A1(_2650_),
    .A2(_2651_),
    .ZN(_2652_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3204_ (.A1(_2650_),
    .A2(_2651_),
    .Z(_2653_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3205_ (.A1(\hvsync_gen.vpos[1] ),
    .A2(_2652_),
    .B(_2590_),
    .ZN(_2654_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3206_ (.A1(_2577_),
    .A2(net107),
    .A3(_2653_),
    .ZN(_2655_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3207_ (.A1(_2654_),
    .A2(_2655_),
    .ZN(_2656_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3208_ (.A1(_2640_),
    .A2(_2656_),
    .Z(_2657_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3209_ (.A1(_2640_),
    .A2(_2656_),
    .ZN(_2658_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai32_1 _3210_ (.A1(net60),
    .A2(_2657_),
    .A3(_2658_),
    .B1(_2645_),
    .B2(_2647_),
    .ZN(\ppp_y__t[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3211_ (.A1(\ppp_x[2] ),
    .A2(\p_p[2] ),
    .ZN(_2659_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3212_ (.A1(\ppp_x[2] ),
    .A2(\p_p[2] ),
    .Z(_2660_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3213_ (.A1(_2643_),
    .A2(_2646_),
    .ZN(_2661_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3214_ (.A1(_2660_),
    .A2(_2661_),
    .ZN(_2662_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3215_ (.A1(_2660_),
    .A2(_2661_),
    .ZN(_2663_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3216_ (.A1(net60),
    .A2(_2662_),
    .ZN(_2664_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3217_ (.A1(net126),
    .A2(net162),
    .ZN(_2665_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _3218_ (.A1(_2648_),
    .A2(_2650_),
    .Z(_2666_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3219_ (.A1(_2648_),
    .A2(_2650_),
    .B(_2665_),
    .ZN(_2667_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3220_ (.A1(_2648_),
    .A2(_2650_),
    .A3(_2665_),
    .Z(_2668_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _3221_ (.A1(_2667_),
    .A2(_2668_),
    .ZN(_2669_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3222_ (.I(_2669_),
    .ZN(_2670_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3223_ (.A1(\hvsync_gen.vpos[2] ),
    .A2(_2670_),
    .ZN(_2671_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3224_ (.A1(\r[13] ),
    .A2(_2671_),
    .ZN(_2672_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3225_ (.A1(\r[13] ),
    .A2(_2671_),
    .Z(_2673_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or3_1 _3226_ (.A1(_2654_),
    .A2(_2657_),
    .A3(_2673_),
    .Z(_2674_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3227_ (.A1(_2654_),
    .A2(_2657_),
    .B(_2673_),
    .ZN(_2675_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3228_ (.A1(_2674_),
    .A2(_2675_),
    .ZN(_2676_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _3229_ (.A1(_2663_),
    .A2(_2664_),
    .B1(_2676_),
    .B2(net61),
    .ZN(\ppp_y__t[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3230_ (.A1(\ppp_x[3] ),
    .A2(\p_p[3] ),
    .ZN(_2677_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3231_ (.A1(\ppp_x[3] ),
    .A2(\p_p[3] ),
    .Z(_2678_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3232_ (.A1(_2659_),
    .A2(_2662_),
    .ZN(_2679_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3233_ (.A1(_2678_),
    .A2(_2679_),
    .ZN(_2680_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3234_ (.A1(_2678_),
    .A2(_2679_),
    .ZN(_2681_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3235_ (.A1(net61),
    .A2(_2680_),
    .ZN(_2682_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3236_ (.A1(_2672_),
    .A2(_2675_),
    .ZN(_2683_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3237_ (.A1(net122),
    .A2(net160),
    .ZN(_2684_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3238_ (.A1(net126),
    .A2(_2570_),
    .B(_2667_),
    .ZN(_2685_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3239_ (.A1(_2684_),
    .A2(_2685_),
    .ZN(_2686_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3240_ (.A1(_2684_),
    .A2(_2685_),
    .Z(_2687_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3241_ (.A1(net96),
    .A2(net43),
    .ZN(_2688_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3242_ (.A1(\r[14] ),
    .A2(_2688_),
    .ZN(_2689_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3243_ (.A1(\r[14] ),
    .A2(_2688_),
    .Z(_2690_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3244_ (.A1(_2683_),
    .A2(_2690_),
    .ZN(_2691_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3245_ (.A1(_2683_),
    .A2(_2690_),
    .ZN(_2692_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _3246_ (.A1(_2681_),
    .A2(_2682_),
    .B1(_2692_),
    .B2(net61),
    .ZN(\ppp_y__t[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3247_ (.A1(\ppp_x[4] ),
    .A2(\p_p[4] ),
    .ZN(_2693_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3248_ (.A1(\ppp_x[4] ),
    .A2(\p_p[4] ),
    .Z(_2694_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3249_ (.A1(_2677_),
    .A2(_2680_),
    .ZN(_2695_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3250_ (.A1(_2694_),
    .A2(_2695_),
    .ZN(_2696_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3251_ (.A1(_2694_),
    .A2(_2695_),
    .ZN(_2697_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3252_ (.A1(net61),
    .A2(_2696_),
    .ZN(_2698_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3253_ (.A1(net85),
    .A2(net157),
    .ZN(_2699_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3254_ (.A1(net116),
    .A2(_2571_),
    .ZN(_2700_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3255_ (.A1(_2699_),
    .A2(_2700_),
    .ZN(_2701_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3256_ (.A1(_2665_),
    .A2(_2684_),
    .Z(_2702_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _3257_ (.A1(_2550_),
    .A2(\hvsync_gen.hpos[1] ),
    .B(\hvsync_gen.hpos[0] ),
    .C(_2551_),
    .ZN(_2703_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _3258_ (.A1(net130),
    .A2(_2567_),
    .B(_2702_),
    .C(_2703_),
    .ZN(_2704_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3259_ (.A1(_2548_),
    .A2(net160),
    .B(net163),
    .ZN(_2705_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _3260_ (.A1(net122),
    .A2(_2569_),
    .B1(_2705_),
    .B2(net126),
    .ZN(_2706_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _3261_ (.A1(_2666_),
    .A2(_2702_),
    .B1(_2704_),
    .B2(_2706_),
    .ZN(_2707_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _3262_ (.A1(_2701_),
    .A2(_2707_),
    .Z(_2708_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3263_ (.A1(net94),
    .A2(_2708_),
    .ZN(_2709_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3264_ (.A1(\r[15] ),
    .A2(_2709_),
    .Z(_2710_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3265_ (.A1(_2689_),
    .A2(_2691_),
    .ZN(_2711_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3266_ (.A1(_2710_),
    .A2(_2711_),
    .ZN(_2712_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3267_ (.A1(_2710_),
    .A2(_2711_),
    .Z(_2713_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai32_1 _3268_ (.A1(net61),
    .A2(_2712_),
    .A3(_2713_),
    .B1(_2697_),
    .B2(_2698_),
    .ZN(\ppp_y__t[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3269_ (.A1(\p_p[5] ),
    .A2(\ppp_x[5] ),
    .ZN(_2714_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3270_ (.A1(_2693_),
    .A2(_2696_),
    .B(_2714_),
    .ZN(_2715_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3271_ (.A1(_2693_),
    .A2(_2696_),
    .A3(_2714_),
    .ZN(_2716_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3272_ (.A1(net60),
    .A2(_2716_),
    .ZN(_2717_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3273_ (.A1(\r[15] ),
    .A2(_2709_),
    .B(_2713_),
    .ZN(_2718_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3274_ (.A1(net112),
    .A2(_2572_),
    .ZN(_2719_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3275_ (.A1(net88),
    .A2(net155),
    .ZN(_2720_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3276_ (.A1(_2719_),
    .A2(_2720_),
    .ZN(_2721_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3277_ (.A1(_2701_),
    .A2(_2707_),
    .B(_2699_),
    .ZN(_2722_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _3278_ (.A1(_2721_),
    .A2(_2722_),
    .Z(_2723_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3279_ (.A1(net93),
    .A2(_2723_),
    .ZN(_2724_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3280_ (.A1(\r[16] ),
    .A2(_2724_),
    .Z(_2725_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3281_ (.I(_2725_),
    .ZN(_2726_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3282_ (.A1(_2718_),
    .A2(_2726_),
    .ZN(_2727_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3283_ (.A1(_2718_),
    .A2(_2726_),
    .ZN(_2728_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _3284_ (.A1(_2715_),
    .A2(_2717_),
    .B1(_2728_),
    .B2(net60),
    .ZN(\ppp_y__t[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3285_ (.A1(\p_p[5] ),
    .A2(\ppp_x[5] ),
    .B(_2715_),
    .ZN(_2729_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3286_ (.A1(\p_p[6] ),
    .A2(\ppp_x[6] ),
    .ZN(_2730_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3287_ (.A1(_2729_),
    .A2(_2730_),
    .ZN(_2731_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3288_ (.A1(_2729_),
    .A2(_2730_),
    .ZN(_2732_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3289_ (.A1(net60),
    .A2(_2732_),
    .ZN(_2733_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3290_ (.A1(_2721_),
    .A2(_2722_),
    .B(_2719_),
    .ZN(_2734_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3291_ (.A1(net153),
    .A2(_2734_),
    .ZN(_2735_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3292_ (.A1(net92),
    .A2(_2735_),
    .ZN(_2736_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3293_ (.A1(\r[17] ),
    .A2(_2736_),
    .Z(_2737_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3294_ (.I(_2737_),
    .ZN(_2738_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3295_ (.A1(\r[16] ),
    .A2(_2724_),
    .B(_2727_),
    .ZN(_2739_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3296_ (.A1(_2738_),
    .A2(_2739_),
    .ZN(_2740_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3297_ (.A1(_2738_),
    .A2(_2739_),
    .ZN(_2741_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _3298_ (.A1(_2731_),
    .A2(_2733_),
    .B1(_2741_),
    .B2(net60),
    .ZN(\ppp_y__t[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3299_ (.A1(\r[17] ),
    .A2(_2736_),
    .B(_2740_),
    .ZN(_2742_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3300_ (.A1(\r[18] ),
    .A2(_2742_),
    .Z(_2743_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3301_ (.A1(\p_p[6] ),
    .A2(\ppp_x[6] ),
    .B(_2731_),
    .ZN(_2744_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3302_ (.A1(\ppp_x[7] ),
    .A2(\p_p[7] ),
    .A3(_2744_),
    .ZN(_2745_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _3303_ (.I0(_2743_),
    .I1(_2745_),
    .S(net60),
    .Z(\ppp_y__t[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3304_ (.A1(_2573_),
    .A2(_2576_),
    .ZN(_2746_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3305_ (.A1(_2573_),
    .A2(_2575_),
    .A3(_2576_),
    .ZN(_2747_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3306_ (.A1(\hvsync_gen.hpos[1] ),
    .A2(\hvsync_gen.hpos[0] ),
    .ZN(_2748_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _3307_ (.A1(net161),
    .A2(net162),
    .A3(net159),
    .A4(net156),
    .ZN(_2749_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3308_ (.A1(_2748_),
    .A2(_2749_),
    .ZN(_2750_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3309_ (.A1(net154),
    .A2(_2750_),
    .ZN(_2751_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _3310_ (.A1(_2574_),
    .A2(_2748_),
    .A3(_2749_),
    .ZN(_2752_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _3311_ (.A1(_2747_),
    .A2(_2752_),
    .ZN(_2753_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _3312_ (.A1(_2747_),
    .A2(_2752_),
    .Z(_2754_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3313_ (.A1(net93),
    .A2(net94),
    .A3(net92),
    .ZN(_2755_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3314_ (.A1(_2581_),
    .A2(_2755_),
    .ZN(_2756_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3315_ (.A1(\hvsync_gen.vpos[8] ),
    .A2(_2756_),
    .ZN(_2757_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3316_ (.A1(\hvsync_gen.vpos[0] ),
    .A2(\hvsync_gen.vpos[1] ),
    .ZN(_2758_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _3317_ (.A1(\hvsync_gen.vpos[0] ),
    .A2(\hvsync_gen.vpos[1] ),
    .A3(net95),
    .A4(net97),
    .ZN(_2759_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3318_ (.A1(_2583_),
    .A2(_2757_),
    .A3(_2759_),
    .ZN(_2760_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3319_ (.A1(net58),
    .A2(_2760_),
    .ZN(_2761_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3320_ (.A1(frame_counter_frac),
    .A2(_2761_),
    .Z(_2762_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3321_ (.A1(net144),
    .A2(_2762_),
    .Z(_2763_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3322_ (.A1(net136),
    .A2(_2763_),
    .Z(_2764_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3323_ (.A1(net127),
    .A2(net131),
    .A3(_2764_),
    .ZN(_2765_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _3324_ (.A1(net131),
    .A2(net136),
    .A3(_2763_),
    .Z(_2766_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3325_ (.A1(net87),
    .A2(_2765_),
    .ZN(_2767_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _3326_ (.A1(net87),
    .A2(_2548_),
    .ZN(_2768_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3327_ (.A1(_2767_),
    .A2(_2768_),
    .ZN(_2769_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3328_ (.A1(net121),
    .A2(net122),
    .ZN(_2770_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3329_ (.A1(_2765_),
    .A2(_2770_),
    .ZN(_2771_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _3330_ (.A1(net167),
    .A2(_2769_),
    .A3(_2771_),
    .ZN(_0081_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3331_ (.I(_0081_),
    .ZN(_0002_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3332_ (.A1(net123),
    .A2(_2765_),
    .ZN(_2772_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3333_ (.A1(net170),
    .A2(_2772_),
    .ZN(_2773_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3334_ (.I(_2773_),
    .ZN(_0080_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3335_ (.A1(_2549_),
    .A2(_2766_),
    .ZN(_2774_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3336_ (.A1(_2773_),
    .A2(_2774_),
    .ZN(_2775_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3337_ (.A1(net170),
    .A2(_2774_),
    .ZN(_2776_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3338_ (.I(_2776_),
    .ZN(_0079_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3339_ (.A1(_0081_),
    .A2(_2776_),
    .B(_2775_),
    .ZN(_0006_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3340_ (.A1(_2765_),
    .A2(_2770_),
    .B(net88),
    .ZN(_2777_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3341_ (.A1(_2546_),
    .A2(net87),
    .ZN(_2778_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3342_ (.A1(net112),
    .A2(net117),
    .ZN(_2779_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3343_ (.A1(net125),
    .A2(net75),
    .ZN(_2780_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _3344_ (.A1(net123),
    .A2(net127),
    .A3(_2766_),
    .A4(net75),
    .ZN(_2781_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _3345_ (.A1(net172),
    .A2(_2777_),
    .A3(_2781_),
    .Z(_0082_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _3346_ (.A1(_0081_),
    .A2(_2776_),
    .A3(_0082_),
    .Z(_2782_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3347_ (.A1(_2775_),
    .A2(_2782_),
    .ZN(_0005_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3348_ (.A1(_0002_),
    .A2(_2772_),
    .A3(_0082_),
    .ZN(_2783_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3349_ (.A1(_0079_),
    .A2(_2783_),
    .ZN(_0007_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3350_ (.A1(_2773_),
    .A2(_2776_),
    .B(_2782_),
    .ZN(_0008_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3351_ (.I(_0008_),
    .ZN(_0009_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3352_ (.A1(_2545_),
    .A2(_2781_),
    .ZN(_2784_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3353_ (.A1(net166),
    .A2(_2784_),
    .ZN(_0083_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3354_ (.A1(_0002_),
    .A2(_0082_),
    .ZN(_2785_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _3355_ (.A1(_0083_),
    .A2(_2785_),
    .Z(_0135_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3356_ (.A1(\frame_counter[7] ),
    .A2(_0082_),
    .Z(_2786_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3357_ (.I(_2786_),
    .ZN(_2787_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3358_ (.A1(_0081_),
    .A2(_2786_),
    .ZN(_0136_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3359_ (.A1(_0135_),
    .A2(_0136_),
    .Z(_0000_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3360_ (.A1(_0081_),
    .A2(_2786_),
    .ZN(_0001_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3361_ (.A1(_0081_),
    .A2(_2786_),
    .ZN(_0003_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3362_ (.A1(_2785_),
    .A2(_2787_),
    .ZN(_0004_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3363_ (.A1(_2597_),
    .A2(_2609_),
    .ZN(_2788_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3364_ (.A1(\r2[1] ),
    .A2(\r1[0] ),
    .ZN(_2789_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _3365_ (.A1(net136),
    .A2(_2788_),
    .A3(_2789_),
    .Z(_2790_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3366_ (.A1(_2788_),
    .A2(_2789_),
    .B(net136),
    .ZN(_2791_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _3367_ (.A1(_2790_),
    .A2(_2791_),
    .Z(\r__t[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3368_ (.A1(net144),
    .A2(_2610_),
    .ZN(_2792_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3369_ (.A1(net144),
    .A2(\r1[1] ),
    .Z(_2793_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3370_ (.A1(\r2[2] ),
    .A2(_2793_),
    .ZN(_2794_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3371_ (.A1(net144),
    .A2(\r2[2] ),
    .A3(\r1[1] ),
    .ZN(_2795_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3372_ (.A1(_2550_),
    .A2(_2795_),
    .ZN(_2796_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3373_ (.A1(_2788_),
    .A2(_2796_),
    .ZN(_2797_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3374_ (.A1(_2788_),
    .A2(_2796_),
    .ZN(_2798_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3375_ (.A1(_2790_),
    .A2(_2798_),
    .ZN(_2799_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _3376_ (.A1(_2790_),
    .A2(_2796_),
    .B1(_2797_),
    .B2(_2799_),
    .ZN(\r__t[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3377_ (.A1(_2788_),
    .A2(_2796_),
    .B(_2799_),
    .ZN(_2800_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3378_ (.A1(net131),
    .A2(_2795_),
    .B(_2794_),
    .ZN(_2801_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3379_ (.A1(net136),
    .A2(_2611_),
    .ZN(_2802_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3380_ (.A1(_2551_),
    .A2(\r1[2] ),
    .ZN(_2803_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3381_ (.A1(net136),
    .A2(\r1[2] ),
    .ZN(_2804_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3382_ (.A1(net137),
    .A2(\r1[2] ),
    .Z(_2805_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3383_ (.A1(net144),
    .A2(_2610_),
    .B(_2805_),
    .ZN(_2806_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3384_ (.A1(_2552_),
    .A2(\r1[1] ),
    .B(_2804_),
    .ZN(_2807_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3385_ (.A1(_2552_),
    .A2(\r1[1] ),
    .A3(_2804_),
    .ZN(_2808_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3386_ (.A1(_2599_),
    .A2(_2806_),
    .A3(_2808_),
    .ZN(_2809_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3387_ (.A1(_2599_),
    .A2(_2792_),
    .A3(_2804_),
    .ZN(_2810_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3388_ (.A1(net127),
    .A2(_2810_),
    .ZN(_2811_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3389_ (.A1(_2801_),
    .A2(_2811_),
    .ZN(_2812_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3390_ (.A1(_2801_),
    .A2(_2811_),
    .ZN(_2813_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3391_ (.A1(_2800_),
    .A2(_2801_),
    .A3(_2811_),
    .ZN(\r__t[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3392_ (.A1(_2549_),
    .A2(_2810_),
    .B(_2809_),
    .ZN(_2814_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3393_ (.A1(net131),
    .A2(_2612_),
    .ZN(_2815_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3394_ (.I(_2815_),
    .ZN(_2816_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3395_ (.A1(net131),
    .A2(\r1[3] ),
    .ZN(_2817_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3396_ (.I(_2817_),
    .ZN(_2818_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3397_ (.A1(_2803_),
    .A2(_2807_),
    .ZN(_2819_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3398_ (.A1(_2803_),
    .A2(_2807_),
    .B(_2818_),
    .ZN(_2820_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3399_ (.A1(_2802_),
    .A2(_2806_),
    .B(_2817_),
    .ZN(_2821_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3400_ (.A1(_2802_),
    .A2(_2806_),
    .A3(_2817_),
    .ZN(_2822_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3401_ (.A1(_2600_),
    .A2(_2820_),
    .A3(_2822_),
    .ZN(_2823_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3402_ (.A1(\r2[4] ),
    .A2(_2818_),
    .A3(_2819_),
    .ZN(_2824_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3403_ (.A1(_2548_),
    .A2(_2824_),
    .ZN(_2825_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3404_ (.A1(_2814_),
    .A2(_2825_),
    .ZN(_2826_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3405_ (.A1(net123),
    .A2(_2814_),
    .A3(_2824_),
    .ZN(_2827_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3406_ (.A1(_2800_),
    .A2(_2813_),
    .B(_2812_),
    .ZN(_2828_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _3407_ (.A1(_2800_),
    .A2(_2813_),
    .B(_2827_),
    .C(_2812_),
    .ZN(_2829_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3408_ (.A1(_2827_),
    .A2(_2828_),
    .ZN(\r__t[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3409_ (.A1(_2826_),
    .A2(_2829_),
    .ZN(_2830_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3410_ (.A1(_2548_),
    .A2(_2824_),
    .B(_2823_),
    .ZN(_2831_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3411_ (.A1(_2549_),
    .A2(\r1[4] ),
    .ZN(_2832_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3412_ (.I(_2832_),
    .ZN(_2833_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3413_ (.A1(net127),
    .A2(\r1[4] ),
    .ZN(_2834_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3414_ (.I(_2834_),
    .ZN(_2835_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3415_ (.A1(_2816_),
    .A2(_2821_),
    .ZN(_2836_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3416_ (.A1(_2816_),
    .A2(_2821_),
    .B(_2835_),
    .ZN(_2837_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3417_ (.A1(_2815_),
    .A2(_2820_),
    .B(_2834_),
    .ZN(_2838_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3418_ (.A1(_2815_),
    .A2(_2820_),
    .A3(_2834_),
    .ZN(_2839_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3419_ (.A1(_2601_),
    .A2(_2837_),
    .A3(_2839_),
    .ZN(_2840_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3420_ (.A1(\r2[5] ),
    .A2(_2835_),
    .A3(_2836_),
    .ZN(_2841_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3421_ (.A1(net87),
    .A2(_2841_),
    .ZN(_2842_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _3422_ (.A1(_2831_),
    .A2(_2842_),
    .Z(_2843_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3423_ (.A1(net87),
    .A2(_2831_),
    .A3(_2841_),
    .ZN(_2844_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3424_ (.A1(_2826_),
    .A2(_2829_),
    .B(_2844_),
    .ZN(_2845_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3425_ (.A1(_2830_),
    .A2(_2844_),
    .ZN(\r__t[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3426_ (.A1(net87),
    .A2(_2841_),
    .B(_2840_),
    .ZN(_2846_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3427_ (.A1(net123),
    .A2(\r1[5] ),
    .ZN(_2847_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3428_ (.A1(net123),
    .A2(\r1[5] ),
    .Z(_2848_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3429_ (.I(_2848_),
    .ZN(_2849_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3430_ (.A1(_2832_),
    .A2(_2838_),
    .ZN(_2850_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3431_ (.A1(_2833_),
    .A2(_2837_),
    .B(_2848_),
    .ZN(_2851_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3432_ (.A1(_2832_),
    .A2(_2838_),
    .A3(_2849_),
    .ZN(_2852_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3433_ (.A1(\r2[6] ),
    .A2(_2851_),
    .A3(_2852_),
    .ZN(_2853_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3434_ (.A1(_2851_),
    .A2(_2852_),
    .B(\r2[6] ),
    .ZN(_2854_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3435_ (.A1(\r2[6] ),
    .A2(_2849_),
    .A3(_2850_),
    .ZN(_2855_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3436_ (.A1(net88),
    .A2(_2855_),
    .ZN(_2856_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3437_ (.A1(_2846_),
    .A2(_2856_),
    .ZN(_2857_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3438_ (.A1(net112),
    .A2(_2846_),
    .A3(_2855_),
    .ZN(_2858_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3439_ (.A1(_2843_),
    .A2(_2845_),
    .B(_2858_),
    .ZN(_2859_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _3440_ (.A1(_2843_),
    .A2(_2845_),
    .A3(_2858_),
    .Z(_2860_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3441_ (.A1(_2859_),
    .A2(_2860_),
    .ZN(\r__t[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3442_ (.A1(_2768_),
    .A2(_2770_),
    .Z(_2861_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3443_ (.A1(_2768_),
    .A2(_2770_),
    .ZN(_2862_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3444_ (.A1(_2614_),
    .A2(net56),
    .ZN(_2863_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3445_ (.A1(\r1[6] ),
    .A2(net57),
    .ZN(_2864_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3446_ (.A1(_2847_),
    .A2(_2851_),
    .ZN(_2865_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3447_ (.A1(_2847_),
    .A2(_2851_),
    .B(_2864_),
    .ZN(_2866_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3448_ (.A1(_2864_),
    .A2(_2865_),
    .ZN(_2867_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3449_ (.A1(\r2[7] ),
    .A2(_2867_),
    .ZN(_2868_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3450_ (.A1(\r2[7] ),
    .A2(_2864_),
    .A3(_2865_),
    .ZN(_2869_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3451_ (.A1(net112),
    .A2(_2854_),
    .B(_2853_),
    .ZN(_2870_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3452_ (.A1(_2869_),
    .A2(_2870_),
    .ZN(_2871_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3453_ (.A1(_2869_),
    .A2(_2870_),
    .Z(_2872_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3454_ (.A1(_2857_),
    .A2(_2859_),
    .ZN(_2873_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3455_ (.A1(_2857_),
    .A2(_2859_),
    .B(_2872_),
    .ZN(_2874_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3456_ (.A1(_2872_),
    .A2(_2873_),
    .ZN(\r__t[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3457_ (.A1(net112),
    .A2(net117),
    .ZN(_2875_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _3458_ (.A1(net112),
    .A2(_2768_),
    .ZN(_2876_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _3459_ (.A1(_2548_),
    .A2(_2875_),
    .ZN(_2877_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3460_ (.A1(net88),
    .A2(_2768_),
    .ZN(_2878_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _3461_ (.I(_2878_),
    .ZN(_2879_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3462_ (.A1(_2615_),
    .A2(_2878_),
    .ZN(_2880_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3463_ (.A1(_2863_),
    .A2(_2866_),
    .ZN(_2881_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3464_ (.A1(_2863_),
    .A2(_2866_),
    .B(_2880_),
    .ZN(_2882_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3465_ (.A1(_2880_),
    .A2(_2881_),
    .ZN(_2883_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3466_ (.A1(\r2[8] ),
    .A2(_2883_),
    .ZN(_2884_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3467_ (.A1(\r2[8] ),
    .A2(_2880_),
    .A3(_2881_),
    .ZN(_2885_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3468_ (.A1(_2868_),
    .A2(_2885_),
    .ZN(_2886_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3469_ (.A1(_2868_),
    .A2(_2885_),
    .ZN(_2887_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3470_ (.A1(_2871_),
    .A2(_2874_),
    .B(_2887_),
    .ZN(_2888_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _3471_ (.A1(_2871_),
    .A2(_2874_),
    .A3(_2887_),
    .Z(_2889_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3472_ (.A1(_2888_),
    .A2(_2889_),
    .ZN(\r__t[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3473_ (.A1(_2886_),
    .A2(_2888_),
    .ZN(_2890_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3474_ (.A1(_2616_),
    .A2(_2877_),
    .ZN(_2891_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3475_ (.A1(_2615_),
    .A2(_2879_),
    .B(_2882_),
    .ZN(_2892_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3476_ (.A1(_2891_),
    .A2(_2892_),
    .Z(_2893_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3477_ (.A1(\r2[9] ),
    .A2(_2893_),
    .ZN(_2894_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _3478_ (.A1(\r2[9] ),
    .A2(_2891_),
    .A3(_2892_),
    .Z(_2895_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3479_ (.A1(\r2[8] ),
    .A2(_2883_),
    .B(_2895_),
    .ZN(_2896_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3480_ (.A1(_2884_),
    .A2(_2895_),
    .ZN(_2897_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3481_ (.A1(_2886_),
    .A2(_2888_),
    .B(_2897_),
    .ZN(_2898_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3482_ (.A1(_2890_),
    .A2(_2897_),
    .ZN(\r__t[9] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3483_ (.A1(\r1[9] ),
    .A2(_2876_),
    .ZN(_2899_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3484_ (.A1(\r1[9] ),
    .A2(_2877_),
    .Z(_2900_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3485_ (.A1(_2616_),
    .A2(_2876_),
    .B(_2882_),
    .ZN(_2901_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _3486_ (.A1(\r1[8] ),
    .A2(_2877_),
    .B1(_2878_),
    .B2(\r1[7] ),
    .C(_2901_),
    .ZN(_2902_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3487_ (.A1(_2900_),
    .A2(_2902_),
    .Z(_2903_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3488_ (.A1(\r2[10] ),
    .A2(_2903_),
    .ZN(_2904_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3489_ (.A1(_2604_),
    .A2(_2900_),
    .A3(_2902_),
    .ZN(_2905_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3490_ (.A1(_2894_),
    .A2(_2905_),
    .ZN(_2906_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3491_ (.A1(_2894_),
    .A2(_2905_),
    .ZN(_2907_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3492_ (.A1(_2896_),
    .A2(_2898_),
    .B(_2907_),
    .ZN(_2908_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _3493_ (.A1(_2896_),
    .A2(_2898_),
    .A3(_2907_),
    .Z(_2909_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3494_ (.A1(_2908_),
    .A2(_2909_),
    .ZN(\r__t[10] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3495_ (.A1(_2900_),
    .A2(_2902_),
    .B(_2899_),
    .ZN(_2910_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3496_ (.A1(net98),
    .A2(_2910_),
    .ZN(_2911_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3497_ (.A1(net98),
    .A2(_2910_),
    .ZN(_2912_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3498_ (.A1(\r2[11] ),
    .A2(_2912_),
    .ZN(_2913_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _3499_ (.A1(\r2[11] ),
    .A2(\r1[10] ),
    .A3(_2910_),
    .Z(_2914_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3500_ (.A1(\r2[10] ),
    .A2(_2903_),
    .B(_2914_),
    .ZN(_2915_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3501_ (.A1(_2904_),
    .A2(_2914_),
    .ZN(_2916_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3502_ (.A1(_2906_),
    .A2(_2908_),
    .ZN(_2917_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3503_ (.A1(_2906_),
    .A2(_2908_),
    .B(_2916_),
    .ZN(_2918_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3504_ (.A1(_2916_),
    .A2(_2917_),
    .ZN(\r__t[11] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _3505_ (.A1(net98),
    .A2(\r1[11] ),
    .A3(_2910_),
    .ZN(_2919_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3506_ (.A1(\r1[11] ),
    .A2(_2911_),
    .Z(_2920_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _3507_ (.A1(\r2[12] ),
    .A2(_2920_),
    .Z(_2921_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3508_ (.A1(\r2[12] ),
    .A2(\r1[11] ),
    .A3(_2911_),
    .ZN(_2922_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3509_ (.I(_2922_),
    .ZN(_2923_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3510_ (.A1(_2913_),
    .A2(_2923_),
    .ZN(_2924_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3511_ (.A1(_2913_),
    .A2(_2922_),
    .Z(_2925_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3512_ (.A1(_2915_),
    .A2(_2918_),
    .B(_2925_),
    .ZN(_2926_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _3513_ (.A1(_2915_),
    .A2(_2918_),
    .A3(_2925_),
    .Z(_2927_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3514_ (.A1(_2926_),
    .A2(_2927_),
    .ZN(\r__t[12] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3515_ (.A1(_2924_),
    .A2(_2926_),
    .ZN(_2928_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3516_ (.A1(_2617_),
    .A2(_2919_),
    .ZN(_2929_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3517_ (.A1(\r1[12] ),
    .A2(_2919_),
    .ZN(_2930_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3518_ (.A1(_2606_),
    .A2(_2930_),
    .ZN(_2931_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3519_ (.A1(_2606_),
    .A2(_2930_),
    .ZN(_2932_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3520_ (.A1(_2921_),
    .A2(_2932_),
    .Z(_2933_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3521_ (.A1(_2921_),
    .A2(_2928_),
    .A3(_2932_),
    .ZN(\r__t[13] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3522_ (.A1(\r1[12] ),
    .A2(\r1[13] ),
    .ZN(_2934_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3523_ (.A1(_2919_),
    .A2(_2934_),
    .ZN(_2935_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3524_ (.A1(\r1[13] ),
    .A2(_2929_),
    .ZN(_2936_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3525_ (.A1(_2607_),
    .A2(_2935_),
    .A3(_2936_),
    .ZN(_2937_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3526_ (.A1(_2607_),
    .A2(\r1[13] ),
    .A3(_2929_),
    .ZN(_2938_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3527_ (.A1(_2931_),
    .A2(_2938_),
    .ZN(_2939_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai33_1 _3528_ (.A1(\r2[12] ),
    .A2(_2920_),
    .A3(_2932_),
    .B1(_2933_),
    .B2(_2924_),
    .B3(_2926_),
    .ZN(_2940_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3529_ (.A1(_2939_),
    .A2(_2940_),
    .ZN(_2941_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3530_ (.A1(_2939_),
    .A2(net5),
    .Z(\r__t[14] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3531_ (.A1(_2931_),
    .A2(_2938_),
    .B(_2941_),
    .ZN(_2942_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3532_ (.A1(\r1[14] ),
    .A2(_2935_),
    .ZN(_2943_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _3533_ (.A1(\r2[15] ),
    .A2(_2943_),
    .Z(_2944_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3534_ (.A1(\r2[15] ),
    .A2(_2943_),
    .ZN(_2945_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3535_ (.A1(_2944_),
    .A2(_2945_),
    .ZN(_2946_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3536_ (.A1(_2937_),
    .A2(_2946_),
    .ZN(_2947_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3537_ (.A1(_2937_),
    .A2(_2946_),
    .Z(_2948_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3538_ (.I(_2948_),
    .ZN(_2949_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3539_ (.A1(_2942_),
    .A2(_2948_),
    .ZN(\r__t[15] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3540_ (.A1(_2942_),
    .A2(_2949_),
    .B(_2947_),
    .ZN(_2950_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3541_ (.A1(\r1[14] ),
    .A2(\r1[15] ),
    .ZN(_2951_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3542_ (.A1(\r1[14] ),
    .A2(\r1[15] ),
    .ZN(_2952_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _3543_ (.I0(_2952_),
    .I1(\r1[15] ),
    .S(_2935_),
    .Z(_2953_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _3544_ (.A1(\r2[16] ),
    .A2(_2953_),
    .Z(_2954_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3545_ (.A1(\r2[16] ),
    .A2(_2953_),
    .ZN(_2955_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3546_ (.A1(_2954_),
    .A2(_2955_),
    .ZN(_2956_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3547_ (.A1(_2944_),
    .A2(_2956_),
    .Z(_2957_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3548_ (.A1(_2944_),
    .A2(_2956_),
    .ZN(_2958_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3549_ (.I(_2958_),
    .ZN(_2959_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3550_ (.A1(_2950_),
    .A2(_2959_),
    .Z(_2960_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3551_ (.A1(_2950_),
    .A2(_2959_),
    .ZN(_2961_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3552_ (.A1(_2960_),
    .A2(_2961_),
    .ZN(\r__t[16] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3553_ (.A1(_2957_),
    .A2(_2960_),
    .ZN(_2962_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3554_ (.A1(_2934_),
    .A2(_2951_),
    .ZN(_2963_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3555_ (.A1(\r1[14] ),
    .A2(\r1[15] ),
    .A3(_2935_),
    .ZN(_2964_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3556_ (.A1(_2618_),
    .A2(_2964_),
    .Z(_2965_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3557_ (.A1(_2618_),
    .A2(_2964_),
    .ZN(_2966_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3558_ (.A1(\r2[17] ),
    .A2(_2966_),
    .ZN(_2967_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3559_ (.A1(_2954_),
    .A2(_2967_),
    .Z(_2968_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3560_ (.A1(_2954_),
    .A2(_2962_),
    .A3(_2967_),
    .ZN(\r__t[17] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3561_ (.A1(\r1[17] ),
    .A2(_2965_),
    .ZN(_2969_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3562_ (.A1(\r1[17] ),
    .A2(_2965_),
    .B(\r2[18] ),
    .ZN(_2970_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3563_ (.A1(_2969_),
    .A2(_2970_),
    .ZN(_2971_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3564_ (.A1(\r2[18] ),
    .A2(\r1[17] ),
    .A3(_2965_),
    .ZN(_2972_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3565_ (.A1(\r2[17] ),
    .A2(_2966_),
    .B(_2972_),
    .ZN(_2973_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or3_1 _3566_ (.A1(\r2[17] ),
    .A2(_2966_),
    .A3(_2972_),
    .Z(_2974_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3567_ (.A1(_2973_),
    .A2(_2974_),
    .ZN(_2975_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai33_1 _3568_ (.A1(\r2[16] ),
    .A2(_2953_),
    .A3(_2967_),
    .B1(_2968_),
    .B2(_2957_),
    .B3(_2960_),
    .ZN(_2976_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3569_ (.A1(_2975_),
    .A2(net2),
    .Z(\r__t[18] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3570_ (.A1(_2975_),
    .A2(_2976_),
    .B(_2973_),
    .ZN(_2977_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3571_ (.A1(_2971_),
    .A2(_2977_),
    .ZN(\r__t[19] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3572_ (.A1(net106),
    .A2(_2620_),
    .ZN(\pp_x_sq__t[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3573_ (.A1(net104),
    .A2(net105),
    .ZN(_2978_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3574_ (.A1(net104),
    .A2(net105),
    .ZN(_2979_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3575_ (.A1(net106),
    .A2(_2979_),
    .ZN(_2980_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3576_ (.A1(_2978_),
    .A2(_2980_),
    .ZN(\pp_x_sq__t[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3577_ (.A1(net106),
    .A2(\dot[3] ),
    .ZN(_2981_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3578_ (.A1(\dot[2] ),
    .A2(\dot[3] ),
    .ZN(_2982_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3579_ (.A1(net104),
    .A2(_2981_),
    .Z(_2983_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3580_ (.A1(\pp_x_sq__t[2] ),
    .A2(_2983_),
    .ZN(\pp_x_sq__t[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3581_ (.A1(net101),
    .A2(net106),
    .ZN(_2984_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3582_ (.A1(\dot[5] ),
    .A2(net106),
    .ZN(_2985_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _3583_ (.A1(net103),
    .A2(net106),
    .B1(net105),
    .B2(\dot[4] ),
    .ZN(_2986_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3584_ (.A1(\dot[5] ),
    .A2(net105),
    .ZN(_2987_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3585_ (.A1(_2619_),
    .A2(_2621_),
    .A3(_2987_),
    .ZN(_2988_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai32_1 _3586_ (.A1(_2619_),
    .A2(_2621_),
    .A3(_2987_),
    .B1(_2986_),
    .B2(_2982_),
    .ZN(_2989_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3587_ (.A1(net100),
    .A2(net106),
    .A3(net73),
    .ZN(_2990_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3588_ (.A1(_2984_),
    .A2(net73),
    .ZN(_2991_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3589_ (.A1(_2984_),
    .A2(_2987_),
    .Z(_2992_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3590_ (.A1(net100),
    .A2(\dot[1] ),
    .ZN(_2993_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3591_ (.A1(net104),
    .A2(\dot[4] ),
    .ZN(_2994_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3592_ (.A1(_2984_),
    .A2(_2987_),
    .A3(_2994_),
    .ZN(_2995_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3593_ (.A1(_2989_),
    .A2(_2995_),
    .ZN(_2996_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3594_ (.A1(_2989_),
    .A2(_2995_),
    .ZN(_2997_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3595_ (.A1(\dot[3] ),
    .A2(_2994_),
    .Z(_2998_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3596_ (.A1(_2987_),
    .A2(_2998_),
    .ZN(_2999_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3597_ (.A1(_2997_),
    .A2(_2999_),
    .ZN(_3000_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3598_ (.A1(_2986_),
    .A2(_2988_),
    .ZN(_3001_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3599_ (.A1(_2982_),
    .A2(_3001_),
    .ZN(_3002_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3600_ (.I(_3002_),
    .ZN(_3003_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3601_ (.A1(_3000_),
    .A2(_3003_),
    .ZN(_3004_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3602_ (.A1(_3000_),
    .A2(_3002_),
    .ZN(_3005_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3603_ (.A1(_2991_),
    .A2(_3005_),
    .Z(_3006_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3604_ (.A1(_2620_),
    .A2(_2621_),
    .A3(_2981_),
    .ZN(_3007_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _3605_ (.A1(net105),
    .A2(\dot[3] ),
    .B1(\dot[4] ),
    .B2(net106),
    .ZN(_3008_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai32_1 _3606_ (.A1(_2620_),
    .A2(_2621_),
    .A3(_2981_),
    .B1(_3008_),
    .B2(_2979_),
    .ZN(_3009_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3607_ (.A1(_3006_),
    .A2(_3009_),
    .ZN(_3010_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3608_ (.A1(_3006_),
    .A2(net72),
    .ZN(_3011_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3609_ (.A1(_3007_),
    .A2(_3008_),
    .ZN(_3012_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _3610_ (.A1(\dot[0] ),
    .A2(net104),
    .A3(\dot[3] ),
    .A4(\dot[4] ),
    .ZN(_3013_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3611_ (.A1(_3011_),
    .A2(_3013_),
    .Z(\pp_x_sq__t[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3612_ (.A1(_3011_),
    .A2(_3013_),
    .B(_3010_),
    .ZN(_3014_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3613_ (.A1(_2991_),
    .A2(_3005_),
    .B(_3004_),
    .ZN(_3015_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3614_ (.I(_3015_),
    .ZN(_3016_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3615_ (.A1(_2997_),
    .A2(_2999_),
    .B(_2996_),
    .ZN(_3017_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _3616_ (.A1(_2985_),
    .A2(_2993_),
    .B1(_2994_),
    .B2(_2992_),
    .ZN(_3018_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3617_ (.A1(net99),
    .A2(\dot[0] ),
    .ZN(_3019_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3618_ (.A1(net99),
    .A2(net105),
    .ZN(_3020_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3619_ (.A1(_2993_),
    .A2(_3019_),
    .ZN(_3021_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3620_ (.A1(_3018_),
    .A2(_3021_),
    .ZN(_3022_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3621_ (.A1(_3018_),
    .A2(_3021_),
    .ZN(_3023_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3622_ (.A1(_3017_),
    .A2(_3023_),
    .ZN(_3024_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3623_ (.A1(_3017_),
    .A2(_3023_),
    .Z(_3025_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _3624_ (.A1(_2621_),
    .A2(_2982_),
    .B1(_2987_),
    .B2(_2998_),
    .ZN(_3026_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3625_ (.A1(net101),
    .A2(net105),
    .A3(_3026_),
    .ZN(_3027_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3626_ (.A1(_2993_),
    .A2(_3026_),
    .ZN(_3028_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3627_ (.A1(net99),
    .A2(\dot[0] ),
    .A3(_3028_),
    .ZN(_3029_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3628_ (.A1(_3019_),
    .A2(_3028_),
    .ZN(_3030_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3629_ (.A1(_3025_),
    .A2(_3030_),
    .ZN(_3031_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3630_ (.A1(_3025_),
    .A2(_3030_),
    .Z(_3032_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3631_ (.A1(_3015_),
    .A2(_3032_),
    .ZN(_3033_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and4_1 _3632_ (.A1(net101),
    .A2(\dot[0] ),
    .A3(net73),
    .A4(_3033_),
    .Z(_3034_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3633_ (.A1(_2990_),
    .A2(_3033_),
    .ZN(_3035_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3634_ (.A1(_3014_),
    .A2(_3035_),
    .ZN(_3036_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3635_ (.A1(_3014_),
    .A2(_3035_),
    .Z(\pp_x_sq__t[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3636_ (.A1(_3016_),
    .A2(_3032_),
    .B(_3034_),
    .ZN(_3037_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3637_ (.I(_3037_),
    .ZN(_3038_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3638_ (.A1(_3027_),
    .A2(_3029_),
    .ZN(_3039_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3639_ (.A1(_3024_),
    .A2(_3031_),
    .ZN(_3040_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3640_ (.A1(net103),
    .A2(net104),
    .ZN(_3041_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3641_ (.A1(_3021_),
    .A2(_3041_),
    .B(_3022_),
    .ZN(_3042_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3642_ (.I(_3042_),
    .ZN(_3043_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3643_ (.A1(net101),
    .A2(net104),
    .ZN(_3044_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3644_ (.A1(net99),
    .A2(net104),
    .ZN(_3045_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3645_ (.A1(_3020_),
    .A2(_3044_),
    .Z(_3046_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _3646_ (.A1(_2984_),
    .A2(_3020_),
    .B1(_3021_),
    .B2(_3041_),
    .ZN(_3047_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3647_ (.A1(_3046_),
    .A2(_3047_),
    .ZN(_3048_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3648_ (.A1(_2621_),
    .A2(_3048_),
    .ZN(_3049_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3649_ (.A1(_2621_),
    .A2(_3048_),
    .ZN(_3050_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3650_ (.A1(_3042_),
    .A2(_3050_),
    .Z(_3051_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3651_ (.I(_3051_),
    .ZN(_3052_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3652_ (.A1(\dot[3] ),
    .A2(\dot[4] ),
    .ZN(_3053_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3653_ (.A1(_3044_),
    .A2(_3053_),
    .Z(_3054_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3654_ (.A1(net101),
    .A2(\dot[4] ),
    .ZN(_3055_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3655_ (.I(_3055_),
    .ZN(_3056_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3656_ (.A1(_3020_),
    .A2(_3044_),
    .A3(_3053_),
    .ZN(_3057_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3657_ (.A1(_3052_),
    .A2(_3057_),
    .ZN(_3058_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3658_ (.A1(_3051_),
    .A2(_3057_),
    .Z(_3059_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3659_ (.I(_3059_),
    .ZN(_3060_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3660_ (.A1(_3040_),
    .A2(_3059_),
    .Z(_3061_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3661_ (.A1(_3027_),
    .A2(_3029_),
    .B(_3061_),
    .ZN(_3062_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3662_ (.A1(_3039_),
    .A2(_3061_),
    .ZN(_3063_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3663_ (.A1(_3038_),
    .A2(_3063_),
    .ZN(_3064_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3664_ (.A1(_3038_),
    .A2(_3063_),
    .ZN(_3065_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _3665_ (.A1(_3036_),
    .A2(_3037_),
    .A3(_3063_),
    .Z(\pp_x_sq__t[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3666_ (.A1(_3036_),
    .A2(_3065_),
    .B(_3064_),
    .ZN(_3066_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3667_ (.A1(_3040_),
    .A2(_3060_),
    .B(_3062_),
    .ZN(_3067_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _3668_ (.A1(_3020_),
    .A2(_3054_),
    .B1(_3055_),
    .B2(_2982_),
    .ZN(_3068_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3669_ (.I(_3068_),
    .ZN(_3069_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3670_ (.A1(_3043_),
    .A2(_3050_),
    .B(_3058_),
    .ZN(_3070_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3671_ (.A1(net103),
    .A2(net100),
    .ZN(_3071_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3672_ (.A1(net103),
    .A2(net100),
    .Z(_3072_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3673_ (.A1(\dot[3] ),
    .A2(_3072_),
    .ZN(_3073_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3674_ (.A1(_3045_),
    .A2(_3073_),
    .ZN(_3074_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3675_ (.A1(_3045_),
    .A2(_3073_),
    .Z(_3075_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3676_ (.A1(_3046_),
    .A2(_3047_),
    .B(_3049_),
    .ZN(_3076_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3677_ (.A1(net99),
    .A2(net104),
    .A3(_2993_),
    .ZN(_3077_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3678_ (.A1(net100),
    .A2(\dot[3] ),
    .ZN(_3078_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3679_ (.I(_3078_),
    .ZN(_3079_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3680_ (.A1(_3077_),
    .A2(_3079_),
    .ZN(_3080_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3681_ (.I(_3080_),
    .ZN(_3081_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3682_ (.A1(_3076_),
    .A2(_3081_),
    .ZN(_0137_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3683_ (.A1(_3076_),
    .A2(_3080_),
    .ZN(_0138_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3684_ (.A1(_3075_),
    .A2(_0138_),
    .Z(_0139_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3685_ (.A1(_3070_),
    .A2(_0139_),
    .ZN(_0140_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3686_ (.A1(_3070_),
    .A2(_0139_),
    .ZN(_0141_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3687_ (.A1(_3069_),
    .A2(_0141_),
    .ZN(_0142_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3688_ (.A1(_3067_),
    .A2(_0142_),
    .Z(_0143_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3689_ (.A1(_3066_),
    .A2(_0143_),
    .ZN(_0144_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3690_ (.A1(_3066_),
    .A2(_0143_),
    .Z(\pp_x_sq__t[9] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3691_ (.A1(_3067_),
    .A2(_0142_),
    .B(_0144_),
    .ZN(_0145_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3692_ (.A1(_3069_),
    .A2(_0141_),
    .B(_0140_),
    .ZN(_0146_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3693_ (.A1(net103),
    .A2(_3079_),
    .B(_3074_),
    .ZN(_0147_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3694_ (.A1(_3075_),
    .A2(_0138_),
    .B(_0137_),
    .ZN(_0148_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3695_ (.I(_0148_),
    .ZN(_0149_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3696_ (.A1(net99),
    .A2(\dot[3] ),
    .ZN(_0150_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3697_ (.A1(_3055_),
    .A2(_0150_),
    .Z(_0151_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3698_ (.A1(net103),
    .A2(_0151_),
    .ZN(_0152_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3699_ (.A1(_2593_),
    .A2(_0151_),
    .ZN(_0153_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3700_ (.A1(_2993_),
    .A2(_3078_),
    .B(_3045_),
    .ZN(_0154_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3701_ (.A1(_0153_),
    .A2(_0154_),
    .ZN(_0155_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3702_ (.I(_0155_),
    .ZN(_0156_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3703_ (.A1(net99),
    .A2(\dot[4] ),
    .ZN(_0157_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3704_ (.A1(_3073_),
    .A2(_0157_),
    .ZN(_0158_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _3705_ (.A1(\dot[7] ),
    .A2(\dot[3] ),
    .B1(\dot[4] ),
    .B2(_3072_),
    .ZN(_0159_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3706_ (.A1(_0158_),
    .A2(_0159_),
    .ZN(_0160_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3707_ (.A1(_0156_),
    .A2(_0160_),
    .ZN(_0161_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3708_ (.A1(_0155_),
    .A2(_0160_),
    .ZN(_0162_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3709_ (.A1(_0149_),
    .A2(_0162_),
    .ZN(_0163_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3710_ (.A1(_0148_),
    .A2(_0162_),
    .ZN(_0164_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3711_ (.I(_0164_),
    .ZN(_0165_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3712_ (.A1(_0147_),
    .A2(_0164_),
    .Z(_0166_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3713_ (.I(_0166_),
    .ZN(_0167_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3714_ (.A1(_0146_),
    .A2(_0167_),
    .ZN(_0168_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3715_ (.A1(_0146_),
    .A2(_0166_),
    .ZN(_0169_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3716_ (.A1(_0145_),
    .A2(_0169_),
    .ZN(_0170_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3717_ (.A1(_0145_),
    .A2(_0169_),
    .Z(\pp_x_sq__t[10] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3718_ (.A1(_0147_),
    .A2(_0165_),
    .B(_0163_),
    .ZN(_0171_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3719_ (.A1(net103),
    .A2(_3056_),
    .B(_0158_),
    .ZN(_0172_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3720_ (.A1(_2593_),
    .A2(\dot[4] ),
    .A3(_0150_),
    .ZN(_0173_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3721_ (.A1(_0153_),
    .A2(_0154_),
    .B(_0173_),
    .ZN(_0174_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _3722_ (.A1(_0156_),
    .A2(_0173_),
    .B1(_0174_),
    .B2(_0161_),
    .ZN(_0175_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3723_ (.A1(_0171_),
    .A2(_0175_),
    .ZN(_0176_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3724_ (.A1(_0171_),
    .A2(_0175_),
    .Z(_0177_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3725_ (.A1(_0168_),
    .A2(_0170_),
    .ZN(_0178_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3726_ (.A1(_0177_),
    .A2(_0178_),
    .ZN(_0179_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3727_ (.A1(_0177_),
    .A2(_0178_),
    .Z(\pp_x_sq__t[11] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3728_ (.A1(_0176_),
    .A2(_0179_),
    .ZN(_0180_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3729_ (.A1(_0152_),
    .A2(_0172_),
    .ZN(_0181_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3730_ (.A1(_3071_),
    .A2(_0157_),
    .B(_0181_),
    .ZN(_0182_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3731_ (.A1(net100),
    .A2(_0182_),
    .ZN(_0183_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _3732_ (.A1(_3071_),
    .A2(_0157_),
    .B1(_0182_),
    .B2(net100),
    .C(_0183_),
    .ZN(_0184_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3733_ (.I(_0184_),
    .ZN(_0185_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3734_ (.A1(net103),
    .A2(net100),
    .A3(_0181_),
    .ZN(_0186_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3735_ (.A1(_3073_),
    .A2(_0157_),
    .B(_0186_),
    .ZN(_0187_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3736_ (.A1(_0184_),
    .A2(_0187_),
    .Z(_0188_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3737_ (.I(_0188_),
    .ZN(_0189_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3738_ (.A1(_0152_),
    .A2(_0155_),
    .B(_0172_),
    .ZN(_0190_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3739_ (.A1(_0189_),
    .A2(_0190_),
    .ZN(_0191_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3740_ (.A1(_0188_),
    .A2(_0190_),
    .ZN(_0192_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3741_ (.A1(_0180_),
    .A2(_0192_),
    .ZN(_0193_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3742_ (.A1(_0180_),
    .A2(_0192_),
    .Z(\pp_x_sq__t[12] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3743_ (.A1(net103),
    .A2(net99),
    .A3(_3055_),
    .ZN(_0194_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _3744_ (.A1(net100),
    .A2(_0182_),
    .B1(_0185_),
    .B2(_0187_),
    .ZN(_0195_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3745_ (.A1(_0194_),
    .A2(_0195_),
    .ZN(_0196_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3746_ (.A1(_0191_),
    .A2(_0193_),
    .B(_0196_),
    .ZN(_0197_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _3747_ (.A1(_0191_),
    .A2(_0193_),
    .A3(_0196_),
    .Z(_0198_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3748_ (.A1(_0197_),
    .A2(_0198_),
    .ZN(\pp_x_sq__t[13] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3749_ (.A1(_2593_),
    .A2(net100),
    .B(_2595_),
    .ZN(_0199_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _3750_ (.I0(_0199_),
    .I1(net102),
    .S(_0197_),
    .Z(\pp_x_sq__t[14] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _3751_ (.I0(_0197_),
    .I1(net99),
    .S(net102),
    .Z(\pp_x_sq__t[15] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3752_ (.A1(net104),
    .A2(net105),
    .A3(_2981_),
    .ZN(_0200_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _3753_ (.A1(_2619_),
    .A2(net105),
    .A3(_2982_),
    .B(_0200_),
    .ZN(_0201_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3754_ (.A1(_3012_),
    .A2(_0201_),
    .Z(\pp_x_sq__t[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3755_ (.A1(_2548_),
    .A2(net126),
    .ZN(_0202_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3756_ (.A1(net122),
    .A2(_2549_),
    .ZN(_0203_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3757_ (.A1(_2634_),
    .A2(_0202_),
    .ZN(_0204_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3758_ (.A1(frame_counter_frac),
    .A2(_2634_),
    .A3(_0202_),
    .ZN(_0205_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3759_ (.A1(_2637_),
    .A2(_0202_),
    .ZN(_0206_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3760_ (.A1(frame_counter_frac),
    .A2(_0206_),
    .B(_0205_),
    .ZN(_0207_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3761_ (.A1(frame_counter_frac),
    .A2(_0206_),
    .B(_2566_),
    .ZN(_0208_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3762_ (.A1(_2566_),
    .A2(_0207_),
    .ZN(_0209_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _3763_ (.A1(\hvsync_gen.vpos[0] ),
    .A2(_0205_),
    .B1(_0209_),
    .B2(net151),
    .ZN(_0210_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3764_ (.A1(net143),
    .A2(_2634_),
    .A3(_0202_),
    .ZN(_0211_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3765_ (.A1(_2638_),
    .A2(_0203_),
    .B(_2552_),
    .ZN(_0212_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3766_ (.A1(_2635_),
    .A2(_0203_),
    .B(net151),
    .ZN(_0213_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3767_ (.A1(_0212_),
    .A2(_0213_),
    .ZN(_0214_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3768_ (.A1(\hvsync_gen.vpos[1] ),
    .A2(_0212_),
    .A3(_0213_),
    .ZN(_0215_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _3769_ (.A1(net143),
    .A2(_0206_),
    .B(_0211_),
    .C(_2577_),
    .ZN(_0216_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3770_ (.A1(_0208_),
    .A2(_0215_),
    .A3(_0216_),
    .ZN(_0217_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3771_ (.A1(_2577_),
    .A2(_0208_),
    .A3(_0214_),
    .ZN(_0218_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3772_ (.A1(_2551_),
    .A2(_0218_),
    .ZN(_0219_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3773_ (.A1(_0210_),
    .A2(_0219_),
    .Z(_0220_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3774_ (.A1(_0210_),
    .A2(_0219_),
    .ZN(_0221_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _3775_ (.A1(_0210_),
    .A2(_0219_),
    .Z(_0222_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3776_ (.A1(_0210_),
    .A2(_0219_),
    .ZN(_0223_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3777_ (.A1(_2544_),
    .A2(_2545_),
    .ZN(_0224_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3778_ (.A1(\frame_counter[8] ),
    .A2(\frame_counter[7] ),
    .ZN(_0225_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3779_ (.A1(_2636_),
    .A2(_0225_),
    .Z(_0226_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3780_ (.A1(_2636_),
    .A2(_0225_),
    .ZN(_0227_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3781_ (.A1(_0222_),
    .A2(net55),
    .ZN(_0228_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3782_ (.A1(_2652_),
    .A2(net55),
    .ZN(_0229_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _3783_ (.A1(net143),
    .A2(_2566_),
    .A3(_0207_),
    .ZN(_0230_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3784_ (.A1(net151),
    .A2(_0209_),
    .ZN(_0231_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3785_ (.A1(net55),
    .A2(_0230_),
    .ZN(_0232_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3786_ (.A1(\frame_counter[8] ),
    .A2(\frame_counter[7] ),
    .ZN(_0233_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3787_ (.A1(_2544_),
    .A2(_2545_),
    .ZN(_0234_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3788_ (.A1(_2630_),
    .A2(_0230_),
    .ZN(_0235_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3789_ (.A1(_2631_),
    .A2(net26),
    .ZN(_0236_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3790_ (.A1(_0235_),
    .A2(_0236_),
    .ZN(_0237_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3791_ (.A1(net87),
    .A2(_0233_),
    .A3(_0237_),
    .ZN(_0238_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3792_ (.A1(_0232_),
    .A2(_0238_),
    .Z(_0239_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3793_ (.A1(_0228_),
    .A2(_0239_),
    .ZN(_0240_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3794_ (.A1(_0228_),
    .A2(_0239_),
    .Z(_0241_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3795_ (.A1(_0229_),
    .A2(_0241_),
    .Z(_0242_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3796_ (.A1(_0222_),
    .A2(net55),
    .A3(_0242_),
    .ZN(_0243_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3797_ (.A1(_0229_),
    .A2(_0239_),
    .ZN(\p_p__t[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3798_ (.A1(_0229_),
    .A2(_0241_),
    .B(_0240_),
    .ZN(_0244_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3799_ (.A1(_2670_),
    .A2(net55),
    .ZN(_0245_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _3800_ (.A1(net118),
    .A2(net71),
    .A3(_0235_),
    .B(_0232_),
    .ZN(_0246_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3801_ (.I(_0246_),
    .ZN(_0247_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3802_ (.A1(net74),
    .A2(_2875_),
    .ZN(_0248_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _3803_ (.A1(net74),
    .A2(_2875_),
    .Z(_0249_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3804_ (.A1(net26),
    .A2(_0249_),
    .ZN(_0250_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3805_ (.A1(_0230_),
    .A2(net54),
    .ZN(_0251_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3806_ (.A1(net87),
    .A2(_0222_),
    .B(_0250_),
    .ZN(_0252_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3807_ (.A1(net118),
    .A2(_0223_),
    .A3(_0251_),
    .ZN(_0253_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3808_ (.A1(_2547_),
    .A2(_0222_),
    .A3(_0250_),
    .ZN(_0254_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3809_ (.A1(net71),
    .A2(_0252_),
    .A3(_0253_),
    .ZN(_0255_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _3810_ (.A1(_2547_),
    .A2(_2652_),
    .B1(net54),
    .B2(net81),
    .ZN(_0256_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _3811_ (.A1(net88),
    .A2(net118),
    .A3(_2630_),
    .A4(_2653_),
    .ZN(_0257_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3812_ (.A1(net70),
    .A2(_0256_),
    .A3(_0257_),
    .ZN(_0258_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _3813_ (.A1(net71),
    .A2(_0252_),
    .A3(_0253_),
    .B(_0258_),
    .ZN(_0259_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3814_ (.I(_0259_),
    .ZN(_0260_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3815_ (.A1(_0255_),
    .A2(_0258_),
    .ZN(_0261_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3816_ (.A1(_0246_),
    .A2(_0261_),
    .ZN(_0262_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3817_ (.A1(_0245_),
    .A2(_0262_),
    .ZN(_0263_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3818_ (.A1(_0245_),
    .A2(_0262_),
    .ZN(_0264_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3819_ (.A1(_0244_),
    .A2(_0264_),
    .ZN(_0265_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3820_ (.A1(_0244_),
    .A2(_0264_),
    .ZN(_0266_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3821_ (.A1(_0243_),
    .A2(_0266_),
    .ZN(_0267_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3822_ (.A1(_0243_),
    .A2(_0266_),
    .Z(\p_p__t[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3823_ (.A1(_0265_),
    .A2(_0267_),
    .ZN(_0268_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3824_ (.A1(_0247_),
    .A2(_0261_),
    .B(_0263_),
    .ZN(_0269_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3825_ (.A1(net43),
    .A2(net55),
    .ZN(_0270_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3826_ (.A1(net137),
    .A2(_0218_),
    .B(_0217_),
    .ZN(_0271_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _3827_ (.I0(_0204_),
    .I1(_0206_),
    .S(_2551_),
    .Z(_0272_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3828_ (.A1(_2578_),
    .A2(_0272_),
    .ZN(_0273_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3829_ (.A1(_2578_),
    .A2(_0272_),
    .ZN(_0274_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3830_ (.A1(_0215_),
    .A2(_0274_),
    .ZN(_0275_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3831_ (.A1(_2578_),
    .A2(_0215_),
    .A3(_0272_),
    .ZN(_0276_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3832_ (.A1(net135),
    .A2(_0276_),
    .ZN(_0277_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3833_ (.A1(_0271_),
    .A2(_0277_),
    .Z(_0278_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3834_ (.A1(_0271_),
    .A2(_0277_),
    .ZN(_0279_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3835_ (.A1(_0271_),
    .A2(_0277_),
    .ZN(_0280_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3836_ (.A1(_0271_),
    .A2(_0277_),
    .Z(_0281_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3837_ (.A1(_0221_),
    .A2(_0281_),
    .ZN(_0282_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3838_ (.A1(_0220_),
    .A2(_0281_),
    .ZN(_0283_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3839_ (.A1(_0227_),
    .A2(_0283_),
    .ZN(_0284_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3840_ (.A1(_0249_),
    .A2(_0283_),
    .ZN(_0285_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3841_ (.A1(net86),
    .A2(_0282_),
    .ZN(_0286_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3842_ (.A1(_0222_),
    .A2(net54),
    .ZN(_0287_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3843_ (.A1(_0286_),
    .A2(_0287_),
    .ZN(_0288_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3844_ (.A1(_0286_),
    .A2(_0287_),
    .ZN(_0289_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _3845_ (.A1(_2779_),
    .A2(net26),
    .B(_0254_),
    .C(_0289_),
    .ZN(_0290_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or4_1 _3846_ (.A1(net118),
    .A2(_0223_),
    .A3(_0251_),
    .A4(_0289_),
    .Z(_0291_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3847_ (.A1(_0233_),
    .A2(_0290_),
    .A3(_0291_),
    .ZN(_0292_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3848_ (.A1(net81),
    .A2(net75),
    .B1(net54),
    .B2(_2652_),
    .ZN(_0293_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3849_ (.A1(net117),
    .A2(_2669_),
    .ZN(_0294_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3850_ (.A1(net117),
    .A2(_2669_),
    .A3(_0293_),
    .ZN(_0295_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3851_ (.A1(_0293_),
    .A2(_0294_),
    .Z(_0296_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3852_ (.I(_0296_),
    .ZN(_0297_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3853_ (.A1(_0257_),
    .A2(_0297_),
    .ZN(_0298_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3854_ (.A1(_0257_),
    .A2(_0297_),
    .B(net80),
    .ZN(_0299_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3855_ (.A1(_0257_),
    .A2(_0297_),
    .B(_0299_),
    .ZN(_0300_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3856_ (.A1(_0292_),
    .A2(_0300_),
    .ZN(_0301_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3857_ (.A1(_0292_),
    .A2(_0300_),
    .Z(_0302_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3858_ (.A1(_0284_),
    .A2(_0302_),
    .Z(_0303_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3859_ (.A1(_0284_),
    .A2(_0292_),
    .A3(_0300_),
    .ZN(_0304_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3860_ (.A1(_0260_),
    .A2(_0304_),
    .ZN(_0305_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3861_ (.A1(_0260_),
    .A2(_0304_),
    .ZN(_0306_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3862_ (.A1(_0259_),
    .A2(_0270_),
    .A3(_0304_),
    .ZN(_0307_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3863_ (.A1(_0269_),
    .A2(_0307_),
    .ZN(_0308_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3864_ (.A1(_0269_),
    .A2(_0307_),
    .ZN(_0309_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3865_ (.A1(_0268_),
    .A2(_0309_),
    .Z(\p_p__t[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3866_ (.A1(_0268_),
    .A2(_0309_),
    .B(_0308_),
    .ZN(_0310_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3867_ (.A1(_0270_),
    .A2(_0306_),
    .B(_0305_),
    .ZN(_0311_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3868_ (.A1(_2708_),
    .A2(_0226_),
    .Z(_0312_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3869_ (.A1(_0284_),
    .A2(_0302_),
    .B(_0301_),
    .ZN(_0313_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3870_ (.A1(_0220_),
    .A2(_0281_),
    .B(_0278_),
    .ZN(_0314_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3871_ (.A1(_0221_),
    .A2(_0280_),
    .B(_0279_),
    .ZN(_0315_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3872_ (.A1(_2550_),
    .A2(_0276_),
    .B(_0275_),
    .ZN(_0316_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3873_ (.A1(net135),
    .A2(_0206_),
    .ZN(_0317_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _3874_ (.A1(net135),
    .A2(_2635_),
    .A3(_0203_),
    .ZN(_0318_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3875_ (.A1(_2550_),
    .A2(_2634_),
    .A3(_0202_),
    .ZN(_0319_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3876_ (.A1(net96),
    .A2(_0318_),
    .Z(_0320_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3877_ (.A1(net96),
    .A2(_0318_),
    .ZN(_0321_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3878_ (.A1(_0320_),
    .A2(_0321_),
    .ZN(_0322_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3879_ (.A1(_0273_),
    .A2(_0317_),
    .A3(_0322_),
    .ZN(_0323_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3880_ (.A1(net126),
    .A2(_0323_),
    .ZN(_0324_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3881_ (.A1(_0316_),
    .A2(_0324_),
    .ZN(_0325_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _3882_ (.A1(_0316_),
    .A2(_0324_),
    .Z(_0326_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3883_ (.A1(_0316_),
    .A2(_0324_),
    .Z(_0327_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3884_ (.A1(_0316_),
    .A2(_0324_),
    .Z(_0328_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3885_ (.A1(_0314_),
    .A2(net17),
    .ZN(_0329_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3886_ (.A1(_0315_),
    .A2(net17),
    .ZN(_0330_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3887_ (.A1(_0226_),
    .A2(_0329_),
    .ZN(_0331_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3888_ (.A1(net54),
    .A2(_0329_),
    .ZN(_0332_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3889_ (.A1(net86),
    .A2(_0285_),
    .A3(_0329_),
    .ZN(_0333_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _3890_ (.A1(_0249_),
    .A2(_0283_),
    .B1(_0330_),
    .B2(net116),
    .ZN(_0334_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _3891_ (.A1(net74),
    .A2(_0222_),
    .B1(_0333_),
    .B2(_0334_),
    .ZN(_0335_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _3892_ (.A1(net85),
    .A2(_0222_),
    .A3(_0285_),
    .A4(_0330_),
    .ZN(_0336_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _3893_ (.A1(net74),
    .A2(_0222_),
    .B1(_0333_),
    .B2(_0334_),
    .C(_0288_),
    .ZN(_0337_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _3894_ (.A1(_0288_),
    .A2(_0291_),
    .A3(_0335_),
    .Z(_0338_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3895_ (.A1(net80),
    .A2(_0338_),
    .Z(_0339_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _3896_ (.A1(net88),
    .A2(net116),
    .A3(_2669_),
    .A4(_2686_),
    .ZN(_0340_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3897_ (.I(_0340_),
    .ZN(_0341_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai222_1 _3898_ (.A1(net116),
    .A2(_2686_),
    .B1(_2779_),
    .B2(_2653_),
    .C1(_0249_),
    .C2(_2669_),
    .ZN(_0342_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3899_ (.A1(_0341_),
    .A2(_0342_),
    .ZN(_0343_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_1 _3900_ (.A1(net116),
    .A2(_2669_),
    .A3(_0293_),
    .A4(_0343_),
    .ZN(_0344_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3901_ (.A1(_0295_),
    .A2(_0343_),
    .Z(_0345_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3902_ (.A1(_0298_),
    .A2(_0345_),
    .ZN(_0346_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3903_ (.A1(_0298_),
    .A2(_0345_),
    .ZN(_0347_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3904_ (.A1(net70),
    .A2(_0347_),
    .ZN(_0348_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3905_ (.A1(_0346_),
    .A2(_0348_),
    .ZN(_0349_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3906_ (.A1(_0339_),
    .A2(_0349_),
    .ZN(_0350_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3907_ (.A1(_0339_),
    .A2(_0349_),
    .ZN(_0351_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3908_ (.A1(_0331_),
    .A2(_0339_),
    .A3(_0349_),
    .ZN(_0352_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3909_ (.A1(_0301_),
    .A2(_0303_),
    .B(_0352_),
    .ZN(_0353_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3910_ (.A1(_0313_),
    .A2(_0352_),
    .Z(_0354_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3911_ (.A1(_0312_),
    .A2(_0313_),
    .A3(_0352_),
    .ZN(_0355_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3912_ (.A1(_0311_),
    .A2(_0355_),
    .ZN(_0356_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3913_ (.A1(_0311_),
    .A2(_0355_),
    .Z(_0357_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3914_ (.A1(_0310_),
    .A2(_0357_),
    .Z(\p_p__t[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3915_ (.A1(_0310_),
    .A2(_0357_),
    .B(_0356_),
    .ZN(_0358_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3916_ (.A1(_0312_),
    .A2(_0354_),
    .B(_0353_),
    .ZN(_0359_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3917_ (.A1(_2723_),
    .A2(_0226_),
    .Z(_0360_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3918_ (.A1(_0331_),
    .A2(_0351_),
    .B(_0350_),
    .ZN(_0361_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3919_ (.A1(_0315_),
    .A2(_0328_),
    .B(_0325_),
    .ZN(_0362_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3920_ (.A1(_0314_),
    .A2(_0327_),
    .B(_0326_),
    .ZN(_0363_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _3921_ (.A1(_2578_),
    .A2(_0272_),
    .B1(_0323_),
    .B2(net126),
    .ZN(_0364_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3922_ (.I(_0364_),
    .ZN(_0365_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3923_ (.A1(net94),
    .A2(_0319_),
    .ZN(_0366_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _3924_ (.A1(_0317_),
    .A2(_0322_),
    .B(_0320_),
    .ZN(_0367_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3925_ (.I(_0367_),
    .ZN(_0368_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3926_ (.A1(net94),
    .A2(_0318_),
    .A3(_0367_),
    .ZN(_0369_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3927_ (.A1(net122),
    .A2(_0369_),
    .Z(_0370_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3928_ (.A1(net122),
    .A2(_0369_),
    .ZN(_0371_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3929_ (.A1(net122),
    .A2(_0369_),
    .ZN(_0372_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3930_ (.A1(_0365_),
    .A2(_0372_),
    .ZN(_0373_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _3931_ (.A1(_0365_),
    .A2(_0372_),
    .Z(_0374_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3932_ (.A1(_0364_),
    .A2(_0372_),
    .ZN(_0375_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3933_ (.A1(_0365_),
    .A2(_0372_),
    .ZN(_0376_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3934_ (.A1(_0362_),
    .A2(_0375_),
    .ZN(_0377_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3935_ (.A1(_0363_),
    .A2(_0375_),
    .ZN(_0378_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3936_ (.A1(_0227_),
    .A2(_0378_),
    .ZN(_0379_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3937_ (.A1(_0291_),
    .A2(_0337_),
    .B(_0336_),
    .ZN(_0380_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3938_ (.A1(net74),
    .A2(_0282_),
    .ZN(_0381_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3939_ (.A1(_0248_),
    .A2(_0377_),
    .ZN(_0382_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3940_ (.A1(net116),
    .A2(_0378_),
    .ZN(_0383_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _3941_ (.A1(net117),
    .A2(_0332_),
    .A3(_0378_),
    .ZN(_0384_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _3942_ (.A1(net54),
    .A2(_0329_),
    .B1(_0377_),
    .B2(net85),
    .ZN(_0385_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3943_ (.A1(_0384_),
    .A2(_0385_),
    .B(_0381_),
    .ZN(_0386_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_1 _3944_ (.A1(net116),
    .A2(_0283_),
    .A3(_0332_),
    .A4(_0377_),
    .ZN(_0387_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _3945_ (.A1(_0384_),
    .A2(_0385_),
    .B(_0333_),
    .C(_0381_),
    .ZN(_0388_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _3946_ (.A1(_0333_),
    .A2(_0380_),
    .A3(_0386_),
    .Z(_0389_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3947_ (.A1(net70),
    .A2(_0389_),
    .ZN(_0390_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _3948_ (.A1(_2669_),
    .A2(_2779_),
    .B1(_0249_),
    .B2(_2686_),
    .ZN(_0391_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3949_ (.A1(net85),
    .A2(_2708_),
    .ZN(_0392_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _3950_ (.A1(net85),
    .A2(_2708_),
    .A3(_0391_),
    .ZN(_0393_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3951_ (.A1(_0391_),
    .A2(_0392_),
    .Z(_0394_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3952_ (.A1(_0340_),
    .A2(_0394_),
    .ZN(_0395_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3953_ (.A1(_0344_),
    .A2(_0347_),
    .A3(_0395_),
    .ZN(_0396_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3954_ (.A1(_0344_),
    .A2(_0347_),
    .B(_0395_),
    .ZN(_0397_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3955_ (.A1(net80),
    .A2(_0397_),
    .ZN(_0398_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _3956_ (.A1(_0396_),
    .A2(_0398_),
    .ZN(_0399_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _3957_ (.A1(net70),
    .A2(_0389_),
    .A3(_0399_),
    .ZN(_0400_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3958_ (.A1(_0390_),
    .A2(_0399_),
    .ZN(_0401_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3959_ (.A1(_0379_),
    .A2(_0401_),
    .ZN(_0402_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3960_ (.A1(_0379_),
    .A2(_0390_),
    .A3(_0399_),
    .ZN(_0403_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3961_ (.A1(_0361_),
    .A2(_0403_),
    .ZN(_0404_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3962_ (.A1(_0361_),
    .A2(_0403_),
    .ZN(_0405_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3963_ (.A1(_0360_),
    .A2(_0361_),
    .A3(_0403_),
    .ZN(_0406_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3964_ (.A1(_0359_),
    .A2(_0406_),
    .ZN(_0407_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3965_ (.A1(_0359_),
    .A2(_0406_),
    .ZN(_0408_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3966_ (.A1(_0358_),
    .A2(_0408_),
    .Z(\p_p__t[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3967_ (.A1(_0358_),
    .A2(_0408_),
    .B(_0407_),
    .ZN(_0409_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3968_ (.A1(_0360_),
    .A2(_0405_),
    .B(_0404_),
    .ZN(_0410_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3969_ (.A1(_2735_),
    .A2(net55),
    .ZN(_0411_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3970_ (.A1(_0379_),
    .A2(_0401_),
    .B(_0400_),
    .ZN(_0412_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _3971_ (.A1(net70),
    .A2(_0389_),
    .A3(_0399_),
    .B(_0402_),
    .ZN(_0413_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3972_ (.A1(net93),
    .A2(_0319_),
    .ZN(_0414_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3973_ (.A1(net93),
    .A2(_0366_),
    .Z(_0415_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _3974_ (.A1(net57),
    .A2(_0415_),
    .Z(_0416_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3975_ (.A1(net57),
    .A2(_0415_),
    .ZN(_0417_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3976_ (.A1(net57),
    .A2(_0415_),
    .ZN(_0418_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3977_ (.A1(_0416_),
    .A2(_0418_),
    .ZN(_0419_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _3978_ (.A1(_0416_),
    .A2(_0418_),
    .B(_0367_),
    .C(_0371_),
    .ZN(_0420_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3979_ (.I(_0420_),
    .ZN(_0421_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _3980_ (.A1(_0367_),
    .A2(_0371_),
    .B(_0416_),
    .C(_0418_),
    .ZN(_0422_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3981_ (.A1(_0368_),
    .A2(_0370_),
    .B(_0419_),
    .ZN(_0423_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3982_ (.A1(_0420_),
    .A2(_0423_),
    .ZN(_0424_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3983_ (.A1(_0362_),
    .A2(_0376_),
    .B(_0374_),
    .ZN(_0425_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3984_ (.A1(_0420_),
    .A2(_0423_),
    .B(_0425_),
    .ZN(_0426_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _3985_ (.A1(_0420_),
    .A2(_0423_),
    .A3(_0425_),
    .Z(_0427_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _3986_ (.A1(_0424_),
    .A2(_0425_),
    .ZN(_0428_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _3987_ (.A1(_0424_),
    .A2(_0425_),
    .Z(_0429_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3988_ (.A1(net55),
    .A2(net12),
    .ZN(_0430_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _3989_ (.A1(_0380_),
    .A2(_0388_),
    .B(_0387_),
    .ZN(_0431_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3990_ (.A1(_0249_),
    .A2(_0429_),
    .ZN(_0432_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _3991_ (.A1(net85),
    .A2(net12),
    .ZN(_0433_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _3992_ (.A1(net54),
    .A2(_0383_),
    .A3(net12),
    .ZN(_0434_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _3993_ (.A1(net117),
    .A2(_0429_),
    .B(_0382_),
    .ZN(_0435_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _3994_ (.A1(net74),
    .A2(_0329_),
    .B1(_0434_),
    .B2(_0435_),
    .ZN(_0436_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_1 _3995_ (.A1(net116),
    .A2(_0330_),
    .A3(_0382_),
    .A4(net12),
    .ZN(_0437_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _3996_ (.I(_0437_),
    .ZN(_0438_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _3997_ (.A1(net74),
    .A2(_0329_),
    .B1(_0434_),
    .B2(_0435_),
    .C(_0384_),
    .ZN(_0439_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _3998_ (.A1(_0384_),
    .A2(_0431_),
    .A3(_0436_),
    .ZN(_0440_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _3999_ (.A1(net70),
    .A2(_0440_),
    .ZN(_0441_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4000_ (.A1(_0341_),
    .A2(_0394_),
    .B(_0397_),
    .ZN(_0442_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _4001_ (.A1(_2687_),
    .A2(net74),
    .B1(net54),
    .B2(_2708_),
    .ZN(_0443_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4002_ (.A1(net85),
    .A2(_2723_),
    .ZN(_0444_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4003_ (.A1(_0443_),
    .A2(_0444_),
    .ZN(_0445_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4004_ (.A1(_0443_),
    .A2(_0444_),
    .ZN(_0446_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4005_ (.A1(_0393_),
    .A2(_0446_),
    .ZN(_0447_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4006_ (.A1(_0393_),
    .A2(_0446_),
    .Z(_0448_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4007_ (.A1(_0442_),
    .A2(_0448_),
    .Z(_0449_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4008_ (.A1(_0442_),
    .A2(_0448_),
    .B(net80),
    .ZN(_0450_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4009_ (.A1(_0449_),
    .A2(_0450_),
    .ZN(_0451_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4010_ (.A1(_0441_),
    .A2(_0451_),
    .Z(_0452_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _4011_ (.A1(_0430_),
    .A2(_0441_),
    .A3(_0451_),
    .Z(_0453_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4012_ (.A1(_0413_),
    .A2(_0453_),
    .Z(_0454_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4013_ (.A1(_0413_),
    .A2(_0453_),
    .Z(_0455_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4014_ (.A1(_0411_),
    .A2(_0412_),
    .A3(_0453_),
    .ZN(_0456_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4015_ (.A1(_0410_),
    .A2(_0456_),
    .Z(_0457_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4016_ (.A1(_0410_),
    .A2(_0456_),
    .Z(_0458_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4017_ (.A1(_0409_),
    .A2(_0458_),
    .Z(\p_p__t[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4018_ (.A1(_0409_),
    .A2(_0458_),
    .B(_0457_),
    .ZN(_0459_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4019_ (.I(_0459_),
    .ZN(_0460_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4020_ (.A1(_0411_),
    .A2(_0455_),
    .B(_0454_),
    .ZN(_0461_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _4021_ (.A1(_2574_),
    .A2(_2734_),
    .B(_2573_),
    .ZN(_0462_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or3_1 _4022_ (.A1(_2573_),
    .A2(_2574_),
    .A3(_2734_),
    .Z(_0463_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4023_ (.A1(_0462_),
    .A2(_0463_),
    .ZN(_0464_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4024_ (.A1(_0462_),
    .A2(_0463_),
    .B(_0227_),
    .ZN(_0465_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai33_1 _4025_ (.A1(net70),
    .A2(_0440_),
    .A3(_0451_),
    .B1(_0452_),
    .B2(_0429_),
    .B3(_0227_),
    .ZN(_0466_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4026_ (.A1(\hvsync_gen.vpos[4] ),
    .A2(_0414_),
    .ZN(_0467_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4027_ (.A1(_0417_),
    .A2(_0467_),
    .ZN(_0468_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4028_ (.A1(net92),
    .A2(_0414_),
    .ZN(_0469_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4029_ (.A1(_2878_),
    .A2(_0469_),
    .ZN(_0470_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4030_ (.A1(_0468_),
    .A2(_0470_),
    .ZN(_0471_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4031_ (.A1(_0468_),
    .A2(_0470_),
    .ZN(_0472_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4032_ (.I(_0472_),
    .ZN(_0473_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _4033_ (.A1(_0363_),
    .A2(_0375_),
    .B(_0422_),
    .C(_0373_),
    .ZN(_0474_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _4034_ (.A1(_0362_),
    .A2(_0376_),
    .B(_0423_),
    .C(_0374_),
    .ZN(_0475_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _4035_ (.A1(_0421_),
    .A2(_0472_),
    .A3(_0474_),
    .ZN(_0476_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4036_ (.A1(_0420_),
    .A2(_0475_),
    .B(_0473_),
    .ZN(_0477_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4037_ (.A1(_0476_),
    .A2(_0477_),
    .Z(_0478_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4038_ (.A1(_0227_),
    .A2(_0478_),
    .ZN(_0479_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4039_ (.A1(_0431_),
    .A2(_0439_),
    .B(_0438_),
    .ZN(_0480_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4040_ (.A1(net116),
    .A2(_0478_),
    .ZN(_0481_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _4041_ (.A1(_0249_),
    .A2(_0433_),
    .A3(_0478_),
    .ZN(_0482_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4042_ (.A1(_0432_),
    .A2(_0481_),
    .ZN(_0483_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4043_ (.A1(_2779_),
    .A2(_0378_),
    .B1(_0482_),
    .B2(_0483_),
    .ZN(_0484_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _4044_ (.A1(_0383_),
    .A2(_0432_),
    .A3(_0484_),
    .Z(_0485_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai221_1 _4045_ (.A1(_2779_),
    .A2(_0378_),
    .B1(_0482_),
    .B2(_0483_),
    .C(_0434_),
    .ZN(_0486_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _4046_ (.A1(_0434_),
    .A2(_0480_),
    .A3(_0484_),
    .Z(_0487_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4047_ (.A1(net70),
    .A2(_0487_),
    .ZN(_0488_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4048_ (.A1(_2708_),
    .A2(net74),
    .B1(net54),
    .B2(_2723_),
    .ZN(_0489_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4049_ (.A1(net85),
    .A2(_2735_),
    .ZN(_0490_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4050_ (.A1(_0489_),
    .A2(_0490_),
    .Z(_0491_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4051_ (.A1(_0489_),
    .A2(_0490_),
    .ZN(_0492_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4052_ (.A1(_0445_),
    .A2(_0492_),
    .ZN(_0493_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _4053_ (.A1(_0447_),
    .A2(_0449_),
    .A3(_0493_),
    .ZN(_0494_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4054_ (.A1(_0447_),
    .A2(_0449_),
    .B(_0493_),
    .ZN(_0495_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4055_ (.A1(net80),
    .A2(_0495_),
    .ZN(_0496_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4056_ (.A1(_0494_),
    .A2(_0496_),
    .ZN(_0497_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _4057_ (.A1(net70),
    .A2(_0487_),
    .A3(_0497_),
    .ZN(_0498_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4058_ (.A1(net70),
    .A2(_0487_),
    .B(_0497_),
    .ZN(_0499_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4059_ (.A1(_0479_),
    .A2(_0488_),
    .A3(_0497_),
    .ZN(_0500_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4060_ (.A1(net3),
    .A2(_0500_),
    .ZN(_0501_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4061_ (.A1(net3),
    .A2(_0500_),
    .ZN(_0502_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _4062_ (.A1(_0465_),
    .A2(_0466_),
    .A3(_0500_),
    .Z(_0503_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4063_ (.A1(_0461_),
    .A2(_0503_),
    .ZN(_0504_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4064_ (.A1(_0461_),
    .A2(_0503_),
    .Z(_0505_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4065_ (.A1(_0459_),
    .A2(_0505_),
    .ZN(\p_p__t[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4066_ (.A1(_0460_),
    .A2(_0505_),
    .B(_0504_),
    .ZN(_0506_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4067_ (.A1(_0465_),
    .A2(_0502_),
    .B(_0501_),
    .ZN(_0507_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4068_ (.A1(_0479_),
    .A2(_0499_),
    .B(_0498_),
    .ZN(_0508_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4069_ (.A1(_0480_),
    .A2(_0486_),
    .B(_0485_),
    .ZN(_0509_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _4070_ (.A1(_0421_),
    .A2(_0472_),
    .A3(_0474_),
    .B(_0471_),
    .ZN(_0510_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4071_ (.A1(net92),
    .A2(_0319_),
    .ZN(_0511_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4072_ (.A1(\hvsync_gen.vpos[5] ),
    .A2(_0511_),
    .ZN(_0512_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4073_ (.A1(_2879_),
    .A2(_0469_),
    .B(_0512_),
    .ZN(_0513_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4074_ (.A1(\hvsync_gen.vpos[7] ),
    .A2(_0511_),
    .ZN(_0514_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4075_ (.A1(_2877_),
    .A2(_0514_),
    .ZN(_0515_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4076_ (.A1(_0513_),
    .A2(_0515_),
    .Z(_0516_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4077_ (.A1(_0513_),
    .A2(_0515_),
    .ZN(_0517_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4078_ (.I(_0517_),
    .ZN(_0518_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _4079_ (.A1(net11),
    .A2(_0517_),
    .ZN(_0519_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4080_ (.A1(net85),
    .A2(_0519_),
    .ZN(_0520_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4081_ (.A1(net88),
    .A2(_0429_),
    .B1(_0478_),
    .B2(_0249_),
    .ZN(_0521_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4082_ (.A1(_0433_),
    .A2(_0521_),
    .ZN(_0522_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4083_ (.A1(_0520_),
    .A2(_0522_),
    .ZN(_0523_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4084_ (.A1(_0509_),
    .A2(_0523_),
    .B(net80),
    .ZN(_0524_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4085_ (.A1(_0509_),
    .A2(_0523_),
    .B(_0524_),
    .ZN(_0525_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _4086_ (.A1(_0443_),
    .A2(_0444_),
    .A3(_0492_),
    .B(_0495_),
    .ZN(_0526_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4087_ (.A1(_2723_),
    .A2(net74),
    .B1(net54),
    .B2(_2735_),
    .ZN(_0527_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4088_ (.A1(net85),
    .A2(_0464_),
    .ZN(_0528_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4089_ (.A1(_0491_),
    .A2(_0528_),
    .Z(_0529_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4090_ (.A1(_0526_),
    .A2(_0527_),
    .A3(_0529_),
    .ZN(_0530_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4091_ (.A1(net80),
    .A2(_0530_),
    .ZN(_0531_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4092_ (.A1(\hvsync_gen.hpos[8] ),
    .A2(_0462_),
    .ZN(_0532_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4093_ (.A1(_2576_),
    .A2(_0462_),
    .ZN(_0533_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4094_ (.A1(net55),
    .A2(_0533_),
    .ZN(_0534_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4095_ (.A1(net55),
    .A2(_0519_),
    .ZN(_0535_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4096_ (.A1(_0531_),
    .A2(_0534_),
    .A3(_0535_),
    .ZN(_0536_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4097_ (.A1(_0525_),
    .A2(_0536_),
    .ZN(_0537_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4098_ (.A1(_0507_),
    .A2(_0508_),
    .A3(_0537_),
    .ZN(_0538_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4099_ (.A1(_0506_),
    .A2(_0538_),
    .Z(\p_p__t[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4100_ (.A1(net141),
    .A2(net149),
    .Z(_0539_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4101_ (.A1(\r[8] ),
    .A2(net78),
    .ZN(_0540_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _4102_ (.A1(net134),
    .A2(net141),
    .A3(net149),
    .Z(_0541_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4103_ (.A1(net141),
    .A2(net149),
    .B(net134),
    .ZN(_0542_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4104_ (.A1(_0541_),
    .A2(_0542_),
    .Z(_0543_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4105_ (.A1(\r[9] ),
    .A2(net69),
    .ZN(_0544_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4106_ (.A1(\r[8] ),
    .A2(net68),
    .ZN(_0545_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4107_ (.A1(\r[9] ),
    .A2(net79),
    .ZN(_0546_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4108_ (.A1(net149),
    .A2(\r[10] ),
    .ZN(_0547_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4109_ (.A1(_0545_),
    .A2(_0546_),
    .Z(_0548_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4110_ (.A1(_0540_),
    .A2(_0544_),
    .B1(_0547_),
    .B2(_0548_),
    .ZN(_0549_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4111_ (.A1(net148),
    .A2(\r[11] ),
    .ZN(_0550_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4112_ (.A1(\r[10] ),
    .A2(net79),
    .ZN(_0551_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4113_ (.A1(_0544_),
    .A2(_0551_),
    .Z(_0552_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4114_ (.A1(\r[10] ),
    .A2(net69),
    .ZN(_0553_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4115_ (.A1(_0544_),
    .A2(_0550_),
    .A3(_0551_),
    .ZN(_0554_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4116_ (.A1(_0549_),
    .A2(_0554_),
    .ZN(_0555_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _4117_ (.A1(net129),
    .A2(net134),
    .A3(net141),
    .A4(net149),
    .ZN(_0556_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4118_ (.A1(_2548_),
    .A2(_0556_),
    .ZN(_0557_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _4119_ (.A1(net87),
    .A2(_2548_),
    .A3(_0556_),
    .ZN(_0558_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4120_ (.A1(net87),
    .A2(_0557_),
    .ZN(_0559_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4121_ (.A1(\r[6] ),
    .A2(net51),
    .ZN(_0560_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4122_ (.A1(_2549_),
    .A2(_0541_),
    .ZN(_0561_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4123_ (.A1(\r[7] ),
    .A2(net66),
    .ZN(_0562_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4124_ (.A1(net125),
    .A2(_0556_),
    .ZN(_0563_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4125_ (.A1(\r[8] ),
    .A2(net64),
    .ZN(_0564_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4126_ (.A1(\r[7] ),
    .A2(net64),
    .ZN(_0565_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4127_ (.A1(\r[8] ),
    .A2(net66),
    .ZN(_0566_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4128_ (.A1(_0565_),
    .A2(_0566_),
    .Z(_0567_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4129_ (.A1(_0560_),
    .A2(_0565_),
    .A3(_0566_),
    .ZN(_0568_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4130_ (.I(_0568_),
    .ZN(_0569_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4131_ (.A1(_0549_),
    .A2(_0554_),
    .ZN(_0570_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4132_ (.A1(_0569_),
    .A2(_0570_),
    .B(_0555_),
    .ZN(_0571_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4133_ (.A1(\r[7] ),
    .A2(net51),
    .ZN(_0572_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4134_ (.A1(\r[9] ),
    .A2(net67),
    .ZN(_0573_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4135_ (.A1(_0564_),
    .A2(_0573_),
    .Z(_0574_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4136_ (.A1(\r[9] ),
    .A2(net64),
    .ZN(_0575_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4137_ (.A1(_0564_),
    .A2(_0572_),
    .A3(_0573_),
    .ZN(_0576_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4138_ (.I(_0576_),
    .ZN(_0577_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4139_ (.A1(_0550_),
    .A2(_0552_),
    .B1(_0553_),
    .B2(_0546_),
    .ZN(_0578_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4140_ (.A1(net148),
    .A2(net107),
    .ZN(_0579_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4141_ (.A1(\r[11] ),
    .A2(net79),
    .ZN(_0580_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4142_ (.A1(\r[11] ),
    .A2(net69),
    .ZN(_0581_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4143_ (.A1(_0553_),
    .A2(_0580_),
    .Z(_0582_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4144_ (.A1(net148),
    .A2(net107),
    .A3(_0582_),
    .ZN(_0583_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4145_ (.A1(_0579_),
    .A2(_0582_),
    .ZN(_0584_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4146_ (.A1(_0578_),
    .A2(_0584_),
    .ZN(_0585_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4147_ (.A1(_0578_),
    .A2(_0584_),
    .ZN(_0586_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4148_ (.A1(_0576_),
    .A2(_0586_),
    .ZN(_0587_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4149_ (.A1(_0571_),
    .A2(_0587_),
    .Z(_0588_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4150_ (.A1(_0562_),
    .A2(_0564_),
    .B1(_0567_),
    .B2(_0560_),
    .ZN(_0589_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _4151_ (.A1(net115),
    .A2(_0558_),
    .ZN(_0590_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4152_ (.A1(_2546_),
    .A2(_0558_),
    .ZN(_0591_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4153_ (.A1(\r[5] ),
    .A2(net50),
    .B1(net48),
    .B2(\r[6] ),
    .ZN(_0592_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4154_ (.I(_0592_),
    .ZN(_0593_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4155_ (.A1(_0589_),
    .A2(_0593_),
    .ZN(_0594_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4156_ (.A1(_0589_),
    .A2(_0592_),
    .ZN(_0595_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4157_ (.A1(_0571_),
    .A2(_0587_),
    .ZN(_0596_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4158_ (.A1(_0588_),
    .A2(_0596_),
    .ZN(_0597_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4159_ (.A1(_0595_),
    .A2(_0597_),
    .B(_0588_),
    .ZN(_0598_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4160_ (.A1(_0572_),
    .A2(_0574_),
    .B1(_0575_),
    .B2(_0566_),
    .ZN(_0599_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4161_ (.A1(\r[6] ),
    .A2(net50),
    .B1(net49),
    .B2(\r[7] ),
    .ZN(_0600_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4162_ (.I(_0600_),
    .ZN(_0601_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4163_ (.A1(_0599_),
    .A2(_0601_),
    .ZN(_0602_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4164_ (.A1(_0599_),
    .A2(_0600_),
    .ZN(_0603_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4165_ (.A1(_0577_),
    .A2(_0586_),
    .B(_0585_),
    .ZN(_0604_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4166_ (.A1(\r[10] ),
    .A2(net65),
    .ZN(_0605_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4167_ (.A1(\r[10] ),
    .A2(net67),
    .ZN(_0606_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4168_ (.A1(_0575_),
    .A2(_0606_),
    .Z(_0607_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4169_ (.A1(\r[8] ),
    .A2(net51),
    .ZN(_0608_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4170_ (.A1(\r[8] ),
    .A2(net51),
    .A3(_0607_),
    .ZN(_0609_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4171_ (.A1(_0607_),
    .A2(_0608_),
    .ZN(_0610_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4172_ (.I(_0610_),
    .ZN(_0611_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4173_ (.A1(_0553_),
    .A2(_0580_),
    .B(_0583_),
    .ZN(_0612_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4174_ (.A1(net107),
    .A2(net69),
    .ZN(_0613_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4175_ (.A1(net107),
    .A2(net79),
    .ZN(_0614_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4176_ (.A1(_0581_),
    .A2(_0614_),
    .Z(_0615_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4177_ (.A1(net150),
    .A2(\r[13] ),
    .ZN(_0616_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4178_ (.A1(_0581_),
    .A2(_0614_),
    .A3(_0616_),
    .ZN(_0617_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4179_ (.A1(_0612_),
    .A2(_0617_),
    .ZN(_0618_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4180_ (.A1(_0612_),
    .A2(_0617_),
    .ZN(_0619_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4181_ (.A1(_0610_),
    .A2(_0619_),
    .ZN(_0620_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4182_ (.A1(_0604_),
    .A2(_0620_),
    .Z(_0621_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4183_ (.A1(_0604_),
    .A2(_0620_),
    .Z(_0622_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4184_ (.A1(_0603_),
    .A2(_0622_),
    .Z(_0623_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4185_ (.I(_0623_),
    .ZN(_0624_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4186_ (.A1(_0598_),
    .A2(_0623_),
    .Z(_0625_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4187_ (.A1(_0594_),
    .A2(_0625_),
    .Z(_0626_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4188_ (.A1(_0598_),
    .A2(_0624_),
    .B(_0626_),
    .ZN(_0627_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4189_ (.A1(_0603_),
    .A2(_0622_),
    .B(_0621_),
    .ZN(_0628_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4190_ (.I(_0628_),
    .ZN(_0629_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4191_ (.A1(_0575_),
    .A2(_0606_),
    .B(_0609_),
    .ZN(_0630_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4192_ (.A1(\r[7] ),
    .A2(_0590_),
    .B1(net48),
    .B2(\r[8] ),
    .ZN(_0631_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4193_ (.I(_0631_),
    .ZN(_0632_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4194_ (.A1(_0630_),
    .A2(_0632_),
    .ZN(_0633_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4195_ (.A1(_0630_),
    .A2(_0631_),
    .ZN(_0634_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4196_ (.A1(_0611_),
    .A2(_0619_),
    .B(_0618_),
    .ZN(_0635_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4197_ (.A1(_0580_),
    .A2(_0613_),
    .B1(_0615_),
    .B2(_0616_),
    .ZN(_0636_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4198_ (.A1(\r[13] ),
    .A2(net69),
    .ZN(_0637_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4199_ (.A1(\r[13] ),
    .A2(net78),
    .ZN(_0638_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4200_ (.A1(_0613_),
    .A2(_0638_),
    .Z(_0639_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4201_ (.A1(net148),
    .A2(\r[14] ),
    .ZN(_0640_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4202_ (.A1(_0613_),
    .A2(_0638_),
    .A3(_0640_),
    .ZN(_0641_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4203_ (.A1(_0636_),
    .A2(_0641_),
    .ZN(_0642_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4204_ (.A1(_0636_),
    .A2(_0641_),
    .ZN(_0643_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4205_ (.A1(\r[11] ),
    .A2(net65),
    .ZN(_0644_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4206_ (.A1(\r[11] ),
    .A2(net67),
    .ZN(_0645_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4207_ (.A1(_0605_),
    .A2(_0645_),
    .Z(_0646_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4208_ (.A1(\r[9] ),
    .A2(net51),
    .ZN(_0647_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4209_ (.A1(_0605_),
    .A2(_0645_),
    .A3(_0647_),
    .ZN(_0648_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4210_ (.I(_0648_),
    .ZN(_0649_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4211_ (.A1(_0643_),
    .A2(_0648_),
    .ZN(_0650_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4212_ (.A1(_0635_),
    .A2(_0650_),
    .Z(_0651_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4213_ (.A1(_0635_),
    .A2(_0650_),
    .ZN(_0652_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4214_ (.A1(_0651_),
    .A2(_0652_),
    .ZN(_0653_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4215_ (.A1(_0634_),
    .A2(_0653_),
    .Z(_0654_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4216_ (.A1(_0629_),
    .A2(_0654_),
    .ZN(_0655_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4217_ (.A1(_0628_),
    .A2(_0654_),
    .Z(_0656_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4218_ (.A1(_0602_),
    .A2(_0656_),
    .Z(_0657_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4219_ (.A1(_0627_),
    .A2(_0657_),
    .ZN(_0658_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4220_ (.A1(_0627_),
    .A2(_0657_),
    .ZN(_0659_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4221_ (.A1(\r[7] ),
    .A2(net78),
    .ZN(_0660_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4222_ (.A1(\r[7] ),
    .A2(net68),
    .ZN(_0661_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4223_ (.A1(net149),
    .A2(\r[9] ),
    .ZN(_0662_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4224_ (.A1(\r[8] ),
    .A2(net78),
    .B1(net68),
    .B2(\r[7] ),
    .ZN(_0663_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4225_ (.A1(_0545_),
    .A2(_0660_),
    .B1(_0662_),
    .B2(_0663_),
    .ZN(_0664_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4226_ (.A1(_0545_),
    .A2(_0546_),
    .A3(_0547_),
    .ZN(_0665_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4227_ (.A1(_0664_),
    .A2(_0665_),
    .ZN(_0666_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4228_ (.A1(\r[5] ),
    .A2(net52),
    .ZN(_0667_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4229_ (.A1(\r[6] ),
    .A2(net66),
    .ZN(_0668_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4230_ (.A1(\r[6] ),
    .A2(net64),
    .ZN(_0669_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4231_ (.A1(_0562_),
    .A2(_0669_),
    .Z(_0670_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4232_ (.A1(_0562_),
    .A2(_0667_),
    .A3(_0669_),
    .ZN(_0671_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4233_ (.A1(_0664_),
    .A2(_0665_),
    .Z(_0672_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4234_ (.A1(_0671_),
    .A2(_0672_),
    .ZN(_0673_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4235_ (.A1(_0666_),
    .A2(_0673_),
    .ZN(_0674_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4236_ (.A1(_0549_),
    .A2(_0554_),
    .A3(_0568_),
    .ZN(_0675_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4237_ (.I(_0675_),
    .ZN(_0676_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4238_ (.A1(_0565_),
    .A2(_0668_),
    .B1(_0670_),
    .B2(_0667_),
    .ZN(_0677_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4239_ (.A1(\r[4] ),
    .A2(net50),
    .B1(net48),
    .B2(\r[5] ),
    .ZN(_0678_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4240_ (.I(_0678_),
    .ZN(_0679_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4241_ (.A1(_0677_),
    .A2(_0679_),
    .ZN(_0680_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4242_ (.A1(_0677_),
    .A2(_0678_),
    .ZN(_0681_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4243_ (.I(_0681_),
    .ZN(_0682_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4244_ (.A1(_0674_),
    .A2(_0676_),
    .ZN(_0683_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4245_ (.A1(_0682_),
    .A2(_0683_),
    .ZN(_0684_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4246_ (.A1(_0674_),
    .A2(_0676_),
    .B(_0684_),
    .ZN(_0685_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4247_ (.I(_0685_),
    .ZN(_0686_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4248_ (.A1(_0595_),
    .A2(_0597_),
    .Z(_0687_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4249_ (.A1(_0686_),
    .A2(_0687_),
    .ZN(_0688_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4250_ (.A1(_0685_),
    .A2(_0687_),
    .Z(_0689_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4251_ (.A1(_0680_),
    .A2(_0689_),
    .Z(_0690_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4252_ (.A1(_0594_),
    .A2(_0625_),
    .ZN(_0691_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4253_ (.A1(_0626_),
    .A2(_0691_),
    .ZN(_0692_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4254_ (.A1(_0688_),
    .A2(_0690_),
    .B(_0692_),
    .ZN(_0693_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4255_ (.A1(_0688_),
    .A2(_0690_),
    .A3(_0692_),
    .ZN(_0694_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4256_ (.I(_0694_),
    .ZN(_0695_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4257_ (.A1(_0680_),
    .A2(_0689_),
    .ZN(_0696_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4258_ (.A1(_0690_),
    .A2(_0696_),
    .ZN(_0697_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4259_ (.A1(\r[6] ),
    .A2(net77),
    .ZN(_0698_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4260_ (.A1(\r[6] ),
    .A2(net68),
    .ZN(_0699_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4261_ (.A1(net149),
    .A2(\r[8] ),
    .ZN(_0700_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4262_ (.A1(\r[7] ),
    .A2(net78),
    .B1(net68),
    .B2(\r[6] ),
    .ZN(_0701_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4263_ (.A1(_0661_),
    .A2(_0698_),
    .B1(_0700_),
    .B2(_0701_),
    .ZN(_0702_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4264_ (.A1(_0540_),
    .A2(_0661_),
    .A3(_0662_),
    .ZN(_0703_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4265_ (.A1(_0702_),
    .A2(_0703_),
    .ZN(_0704_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4266_ (.A1(\r[4] ),
    .A2(net52),
    .ZN(_0705_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4267_ (.A1(\r[5] ),
    .A2(net64),
    .ZN(_0706_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4268_ (.A1(_0668_),
    .A2(_0706_),
    .Z(_0707_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4269_ (.A1(\r[5] ),
    .A2(net66),
    .ZN(_0708_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4270_ (.A1(_0668_),
    .A2(_0705_),
    .A3(_0706_),
    .ZN(_0709_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _4271_ (.A1(_0702_),
    .A2(_0703_),
    .Z(_0710_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4272_ (.A1(_0709_),
    .A2(_0710_),
    .ZN(_0711_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4273_ (.A1(_0704_),
    .A2(_0711_),
    .ZN(_0712_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4274_ (.A1(_0671_),
    .A2(_0672_),
    .Z(_0713_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4275_ (.A1(_0712_),
    .A2(_0713_),
    .Z(_0714_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4276_ (.A1(_0705_),
    .A2(_0707_),
    .B1(_0708_),
    .B2(_0669_),
    .ZN(_0715_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4277_ (.A1(net108),
    .A2(net50),
    .B1(net48),
    .B2(\r[4] ),
    .ZN(_0716_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4278_ (.I(_0716_),
    .ZN(_0717_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4279_ (.A1(_0715_),
    .A2(_0717_),
    .ZN(_0718_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4280_ (.A1(_0715_),
    .A2(_0716_),
    .ZN(_0719_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4281_ (.A1(_0712_),
    .A2(_0713_),
    .Z(_0720_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4282_ (.A1(_0719_),
    .A2(_0720_),
    .B(_0714_),
    .ZN(_0721_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4283_ (.A1(_0682_),
    .A2(_0683_),
    .ZN(_0722_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4284_ (.A1(_0721_),
    .A2(_0722_),
    .ZN(_0723_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4285_ (.A1(_0718_),
    .A2(_0723_),
    .Z(_0724_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4286_ (.A1(_0721_),
    .A2(_0722_),
    .B(_0724_),
    .ZN(_0725_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _4287_ (.A1(_0690_),
    .A2(_0696_),
    .A3(_0725_),
    .Z(_0726_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4288_ (.A1(\r[5] ),
    .A2(net77),
    .ZN(_0727_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4289_ (.A1(\r[5] ),
    .A2(_0541_),
    .A3(_0542_),
    .ZN(_0728_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4290_ (.A1(net149),
    .A2(\r[7] ),
    .ZN(_0729_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4291_ (.A1(_0698_),
    .A2(_0728_),
    .Z(_0730_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4292_ (.A1(_0699_),
    .A2(_0727_),
    .B1(_0729_),
    .B2(_0730_),
    .ZN(_0731_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4293_ (.A1(_0660_),
    .A2(_0699_),
    .A3(_0700_),
    .ZN(_0732_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4294_ (.A1(_0731_),
    .A2(_0732_),
    .ZN(_0733_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4295_ (.A1(_0731_),
    .A2(_0732_),
    .ZN(_0734_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4296_ (.A1(net108),
    .A2(net52),
    .ZN(_0735_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4297_ (.A1(\r[4] ),
    .A2(net66),
    .ZN(_0736_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4298_ (.A1(\r[4] ),
    .A2(net64),
    .ZN(_0737_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4299_ (.A1(_0708_),
    .A2(_0737_),
    .Z(_0738_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4300_ (.A1(net108),
    .A2(net52),
    .A3(_0738_),
    .ZN(_0739_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4301_ (.A1(_0735_),
    .A2(_0738_),
    .Z(_0740_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4302_ (.A1(_0734_),
    .A2(_0740_),
    .B(_0733_),
    .ZN(_0741_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4303_ (.A1(_0709_),
    .A2(_0710_),
    .Z(_0742_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4304_ (.A1(_0741_),
    .A2(_0742_),
    .Z(_0743_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4305_ (.A1(_0708_),
    .A2(_0737_),
    .B(_0739_),
    .ZN(_0744_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4306_ (.A1(net109),
    .A2(net50),
    .B1(net48),
    .B2(net108),
    .ZN(_0745_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4307_ (.I(_0745_),
    .ZN(_0746_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4308_ (.A1(_0744_),
    .A2(_0746_),
    .ZN(_0747_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4309_ (.I(_0747_),
    .ZN(_0748_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4310_ (.A1(_0744_),
    .A2(_0745_),
    .ZN(_0749_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4311_ (.A1(_0741_),
    .A2(_0742_),
    .Z(_0750_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4312_ (.A1(_0749_),
    .A2(_0750_),
    .B(_0743_),
    .ZN(_0751_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4313_ (.A1(_0719_),
    .A2(_0720_),
    .ZN(_0752_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4314_ (.A1(_0751_),
    .A2(_0752_),
    .Z(_0753_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4315_ (.A1(_0748_),
    .A2(_0753_),
    .ZN(_0754_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4316_ (.A1(_0751_),
    .A2(_0752_),
    .B(_0754_),
    .ZN(_0755_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4317_ (.A1(_0718_),
    .A2(_0723_),
    .Z(_0756_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4318_ (.A1(_0755_),
    .A2(_0756_),
    .ZN(_0757_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4319_ (.A1(\r[4] ),
    .A2(net77),
    .ZN(_0758_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4320_ (.A1(\r[4] ),
    .A2(_0541_),
    .A3(_0542_),
    .ZN(_0759_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4321_ (.A1(net149),
    .A2(\r[6] ),
    .ZN(_0760_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4322_ (.A1(_0727_),
    .A2(_0759_),
    .Z(_0761_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4323_ (.A1(_0728_),
    .A2(_0758_),
    .B1(_0760_),
    .B2(_0761_),
    .ZN(_0762_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4324_ (.A1(_0698_),
    .A2(_0728_),
    .A3(_0729_),
    .ZN(_0763_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4325_ (.A1(_0762_),
    .A2(_0763_),
    .ZN(_0764_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4326_ (.A1(_0762_),
    .A2(_0763_),
    .ZN(_0765_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4327_ (.A1(net109),
    .A2(net52),
    .ZN(_0766_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4328_ (.A1(net108),
    .A2(net66),
    .ZN(_0767_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4329_ (.A1(\r[3] ),
    .A2(net64),
    .ZN(_0768_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4330_ (.A1(_0736_),
    .A2(_0768_),
    .Z(_0769_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4331_ (.A1(net109),
    .A2(net52),
    .A3(_0769_),
    .ZN(_0770_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4332_ (.A1(_0766_),
    .A2(_0769_),
    .Z(_0771_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4333_ (.A1(_0765_),
    .A2(_0771_),
    .B(_0764_),
    .ZN(_0772_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4334_ (.A1(_0734_),
    .A2(_0740_),
    .Z(_0773_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4335_ (.A1(_0772_),
    .A2(_0773_),
    .Z(_0774_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4336_ (.A1(_0736_),
    .A2(_0768_),
    .B(_0770_),
    .ZN(_0775_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4337_ (.A1(net110),
    .A2(net50),
    .B1(net48),
    .B2(net109),
    .ZN(_0776_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4338_ (.I(_0776_),
    .ZN(_0777_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4339_ (.A1(_0775_),
    .A2(_0777_),
    .ZN(_0778_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4340_ (.I(_0778_),
    .ZN(_0779_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4341_ (.A1(_0775_),
    .A2(_0776_),
    .ZN(_0780_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4342_ (.A1(_0772_),
    .A2(_0773_),
    .Z(_0781_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4343_ (.A1(_0780_),
    .A2(_0781_),
    .B(_0774_),
    .ZN(_0782_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4344_ (.A1(_0749_),
    .A2(_0750_),
    .ZN(_0783_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4345_ (.A1(_0782_),
    .A2(_0783_),
    .ZN(_0784_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4346_ (.A1(_0782_),
    .A2(_0783_),
    .Z(_0785_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4347_ (.A1(_0779_),
    .A2(_0785_),
    .B(_0784_),
    .ZN(_0786_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4348_ (.A1(_0748_),
    .A2(_0753_),
    .ZN(_0787_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4349_ (.A1(_0786_),
    .A2(_0787_),
    .ZN(_0788_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4350_ (.A1(net108),
    .A2(net77),
    .ZN(_0789_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4351_ (.A1(net108),
    .A2(net68),
    .ZN(_0790_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4352_ (.A1(net147),
    .A2(\r[5] ),
    .ZN(_0791_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4353_ (.A1(\r[4] ),
    .A2(net77),
    .B1(net68),
    .B2(net108),
    .ZN(_0792_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4354_ (.A1(_0759_),
    .A2(_0789_),
    .B1(_0791_),
    .B2(_0792_),
    .ZN(_0793_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4355_ (.A1(_0727_),
    .A2(_0759_),
    .A3(_0760_),
    .ZN(_0794_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4356_ (.A1(_0793_),
    .A2(_0794_),
    .ZN(_0795_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4357_ (.A1(_0793_),
    .A2(_0794_),
    .ZN(_0796_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4358_ (.A1(net110),
    .A2(net52),
    .ZN(_0797_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4359_ (.A1(\r[2] ),
    .A2(net66),
    .ZN(_0798_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4360_ (.A1(net109),
    .A2(net64),
    .ZN(_0799_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4361_ (.A1(_0767_),
    .A2(_0799_),
    .Z(_0800_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4362_ (.A1(net110),
    .A2(net52),
    .A3(_0800_),
    .ZN(_0801_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4363_ (.A1(_0797_),
    .A2(_0800_),
    .Z(_0802_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4364_ (.A1(_0796_),
    .A2(_0802_),
    .B(_0795_),
    .ZN(_0803_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4365_ (.A1(_0765_),
    .A2(_0771_),
    .Z(_0804_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4366_ (.A1(_0803_),
    .A2(_0804_),
    .Z(_0805_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4367_ (.A1(_0767_),
    .A2(_0799_),
    .B(_0801_),
    .ZN(_0806_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4368_ (.A1(net110),
    .A2(net48),
    .ZN(_0807_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4369_ (.A1(\r[0] ),
    .A2(net50),
    .ZN(_0808_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4370_ (.A1(_0807_),
    .A2(_0808_),
    .ZN(_0809_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4371_ (.A1(_0806_),
    .A2(_0809_),
    .ZN(_0810_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4372_ (.I(_0810_),
    .ZN(_0811_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4373_ (.A1(_0806_),
    .A2(_0809_),
    .Z(_0812_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4374_ (.A1(_0803_),
    .A2(_0804_),
    .Z(_0813_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4375_ (.A1(_0812_),
    .A2(_0813_),
    .B(_0805_),
    .ZN(_0814_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4376_ (.A1(_0772_),
    .A2(_0773_),
    .A3(_0780_),
    .ZN(_0815_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4377_ (.A1(_0814_),
    .A2(_0815_),
    .ZN(_0816_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4378_ (.A1(_0814_),
    .A2(_0815_),
    .Z(_0817_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4379_ (.A1(_0811_),
    .A2(_0817_),
    .B(_0816_),
    .ZN(_0818_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4380_ (.A1(_0779_),
    .A2(_0785_),
    .ZN(_0819_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4381_ (.A1(_0818_),
    .A2(_0819_),
    .ZN(_0820_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4382_ (.A1(_0810_),
    .A2(_0817_),
    .ZN(_0821_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4383_ (.A1(net109),
    .A2(net77),
    .ZN(_0822_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4384_ (.A1(net109),
    .A2(net68),
    .ZN(_0823_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4385_ (.A1(net147),
    .A2(\r[4] ),
    .ZN(_0824_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4386_ (.A1(net108),
    .A2(net77),
    .B1(net68),
    .B2(net109),
    .ZN(_0825_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4387_ (.A1(_0790_),
    .A2(_0822_),
    .B1(_0824_),
    .B2(_0825_),
    .ZN(_0826_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4388_ (.A1(_0758_),
    .A2(_0790_),
    .A3(_0791_),
    .ZN(_0827_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4389_ (.A1(_0826_),
    .A2(_0827_),
    .ZN(_0828_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4390_ (.A1(_0826_),
    .A2(_0827_),
    .ZN(_0829_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4391_ (.A1(\r[0] ),
    .A2(net52),
    .ZN(_0830_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4392_ (.A1(\r[1] ),
    .A2(net64),
    .ZN(_0831_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4393_ (.A1(_0798_),
    .A2(_0831_),
    .Z(_0832_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4394_ (.A1(\r[0] ),
    .A2(net52),
    .A3(_0832_),
    .ZN(_0833_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4395_ (.A1(_0830_),
    .A2(_0832_),
    .Z(_0834_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4396_ (.A1(_0829_),
    .A2(_0834_),
    .B(_0828_),
    .ZN(_0835_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4397_ (.A1(_0793_),
    .A2(_0794_),
    .A3(_0802_),
    .ZN(_0836_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4398_ (.A1(_0835_),
    .A2(_0836_),
    .ZN(_0837_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4399_ (.A1(_0798_),
    .A2(_0831_),
    .B(_0833_),
    .ZN(_0838_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4400_ (.A1(\r[0] ),
    .A2(net48),
    .ZN(_0839_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4401_ (.A1(\r[0] ),
    .A2(net48),
    .A3(_0838_),
    .ZN(_0840_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4402_ (.A1(_0838_),
    .A2(_0839_),
    .Z(_0841_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4403_ (.A1(_0835_),
    .A2(_0836_),
    .ZN(_0842_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4404_ (.A1(_0841_),
    .A2(_0842_),
    .B(_0837_),
    .ZN(_0843_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _4405_ (.A1(_0803_),
    .A2(_0804_),
    .A3(_0812_),
    .Z(_0844_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4406_ (.A1(_0843_),
    .A2(_0844_),
    .ZN(_0845_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4407_ (.A1(\r[0] ),
    .A2(net66),
    .ZN(_0846_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4408_ (.A1(_0831_),
    .A2(_0846_),
    .ZN(_0847_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4409_ (.A1(net110),
    .A2(net66),
    .B1(net64),
    .B2(\r[0] ),
    .ZN(_0848_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4410_ (.A1(_0847_),
    .A2(_0848_),
    .Z(_0849_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4411_ (.A1(net110),
    .A2(net77),
    .ZN(_0850_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4412_ (.A1(net110),
    .A2(_0541_),
    .A3(_0542_),
    .ZN(_0851_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4413_ (.A1(net147),
    .A2(net108),
    .ZN(_0852_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4414_ (.A1(_0822_),
    .A2(_0851_),
    .ZN(_0853_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4415_ (.A1(_0823_),
    .A2(_0850_),
    .B1(_0852_),
    .B2(_0853_),
    .ZN(_0854_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4416_ (.A1(_0789_),
    .A2(_0823_),
    .A3(_0824_),
    .ZN(_0855_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4417_ (.A1(_0854_),
    .A2(_0855_),
    .ZN(_0856_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4418_ (.A1(_0854_),
    .A2(_0855_),
    .ZN(_0857_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4419_ (.A1(_0849_),
    .A2(_0857_),
    .Z(_0858_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4420_ (.A1(_0849_),
    .A2(_0857_),
    .ZN(_0859_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4421_ (.A1(_0858_),
    .A2(_0859_),
    .ZN(_0860_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4422_ (.A1(_0852_),
    .A2(_0853_),
    .Z(_0861_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4423_ (.A1(net147),
    .A2(net109),
    .B1(net110),
    .B2(net77),
    .ZN(_0862_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _4424_ (.A1(_2551_),
    .A2(net144),
    .A3(net109),
    .A4(net110),
    .ZN(_0863_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4425_ (.A1(\r[0] ),
    .A2(net68),
    .ZN(_0864_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4426_ (.A1(_0862_),
    .A2(_0864_),
    .B(_0863_),
    .ZN(_0865_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4427_ (.A1(_0861_),
    .A2(_0865_),
    .ZN(_0866_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4428_ (.A1(_0861_),
    .A2(_0865_),
    .Z(_0867_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4429_ (.A1(\r[0] ),
    .A2(net66),
    .A3(_0867_),
    .ZN(_0868_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4430_ (.A1(_0866_),
    .A2(_0868_),
    .Z(_0869_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4431_ (.A1(_0860_),
    .A2(_0869_),
    .ZN(_0870_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _4432_ (.A1(net110),
    .A2(\r[0] ),
    .A3(net77),
    .A4(_0853_),
    .ZN(_0871_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4433_ (.A1(_0846_),
    .A2(_0867_),
    .Z(_0872_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai32_1 _4434_ (.A1(_2552_),
    .A2(_0871_),
    .A3(_0872_),
    .B1(_0860_),
    .B2(_0869_),
    .ZN(_0873_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _4435_ (.A1(_0826_),
    .A2(_0827_),
    .A3(_0834_),
    .Z(_0874_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4436_ (.A1(_0856_),
    .A2(_0858_),
    .A3(_0874_),
    .ZN(_0875_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4437_ (.A1(_0856_),
    .A2(_0858_),
    .B(_0874_),
    .ZN(_0876_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _4438_ (.A1(_0870_),
    .A2(net16),
    .B1(_0875_),
    .B2(_0847_),
    .C(_0876_),
    .ZN(_0877_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4439_ (.A1(_0841_),
    .A2(_0842_),
    .Z(_0878_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4440_ (.A1(_0841_),
    .A2(_0842_),
    .B1(_0847_),
    .B2(_0875_),
    .ZN(_0879_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _4441_ (.A1(_0847_),
    .A2(_0870_),
    .A3(_0873_),
    .A4(_0876_),
    .ZN(_0880_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _4442_ (.A1(_0877_),
    .A2(_0878_),
    .A3(_0879_),
    .B(_0880_),
    .ZN(_0881_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4443_ (.A1(_0843_),
    .A2(_0844_),
    .ZN(_0882_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4444_ (.A1(_0840_),
    .A2(_0882_),
    .B(_0845_),
    .ZN(_0883_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4445_ (.A1(_0821_),
    .A2(_0883_),
    .ZN(_0884_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4446_ (.A1(_0840_),
    .A2(_0843_),
    .A3(_0844_),
    .ZN(_0885_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4447_ (.A1(_0821_),
    .A2(_0883_),
    .B1(_0885_),
    .B2(_0881_),
    .ZN(_0886_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4448_ (.A1(_0884_),
    .A2(_0886_),
    .ZN(_0887_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai32_1 _4449_ (.A1(_0820_),
    .A2(_0884_),
    .A3(_0886_),
    .B1(_0819_),
    .B2(_0818_),
    .ZN(_0888_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4450_ (.A1(_0786_),
    .A2(_0787_),
    .ZN(_0889_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _4451_ (.A1(net10),
    .A2(_0889_),
    .B(_0788_),
    .ZN(_0890_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4452_ (.A1(_0755_),
    .A2(_0756_),
    .ZN(_0891_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _4453_ (.A1(_0890_),
    .A2(_0891_),
    .B(_0757_),
    .ZN(_0892_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4454_ (.A1(_0697_),
    .A2(_0725_),
    .ZN(_0893_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4455_ (.A1(_0892_),
    .A2(_0893_),
    .B(_0726_),
    .ZN(_0894_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _4456_ (.A1(_0892_),
    .A2(_0893_),
    .B(_0693_),
    .C(_0726_),
    .ZN(_0895_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4457_ (.A1(_0695_),
    .A2(_0895_),
    .ZN(_0896_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4458_ (.A1(_0659_),
    .A2(_0896_),
    .Z(_0897_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4459_ (.A1(_0693_),
    .A2(_0695_),
    .ZN(_0898_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4460_ (.A1(_0894_),
    .A2(_0898_),
    .Z(_0899_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _4461_ (.I0(_0897_),
    .I1(_0899_),
    .S(net56),
    .Z(_0900_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _4462_ (.A1(_0786_),
    .A2(_0787_),
    .A3(net9),
    .Z(_0901_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _4463_ (.A1(net121),
    .A2(net125),
    .B(net114),
    .ZN(_0902_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4464_ (.A1(_2546_),
    .A2(_2770_),
    .ZN(_0903_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4465_ (.A1(_0820_),
    .A2(_0887_),
    .ZN(_0904_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4466_ (.A1(net56),
    .A2(_0901_),
    .B1(_0904_),
    .B2(_2768_),
    .ZN(_0905_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _4467_ (.A1(net125),
    .A2(net75),
    .B(_0902_),
    .ZN(_0906_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4468_ (.A1(_2780_),
    .A2(_0903_),
    .ZN(_0907_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _4469_ (.A1(_0755_),
    .A2(_0756_),
    .A3(_0890_),
    .Z(_0908_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4470_ (.A1(net56),
    .A2(_0908_),
    .ZN(_0909_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4471_ (.A1(_0892_),
    .A2(_0893_),
    .Z(_0910_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4472_ (.A1(net56),
    .A2(_0910_),
    .B(_0909_),
    .ZN(_0911_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4473_ (.A1(_2780_),
    .A2(_0900_),
    .B1(_0907_),
    .B2(_0911_),
    .ZN(_0912_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4474_ (.I(_0912_),
    .ZN(_0913_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4475_ (.A1(_0903_),
    .A2(_0905_),
    .B(_0913_),
    .ZN(\dot__t[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _4476_ (.A1(_0659_),
    .A2(_0695_),
    .A3(_0895_),
    .B(_0658_),
    .ZN(_0914_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4477_ (.A1(_0602_),
    .A2(_0656_),
    .B(_0655_),
    .ZN(_0915_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4478_ (.I(_0915_),
    .ZN(_0916_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4479_ (.A1(_0634_),
    .A2(_0653_),
    .B(_0651_),
    .ZN(_0917_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4480_ (.I(_0917_),
    .ZN(_0918_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4481_ (.A1(_0606_),
    .A2(_0644_),
    .B1(_0646_),
    .B2(_0647_),
    .ZN(_0919_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4482_ (.A1(\r[8] ),
    .A2(_0590_),
    .B1(net49),
    .B2(\r[9] ),
    .ZN(_0920_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4483_ (.I(_0920_),
    .ZN(_0921_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4484_ (.A1(_0919_),
    .A2(_0921_),
    .ZN(_0922_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4485_ (.A1(_0919_),
    .A2(_0920_),
    .ZN(_0923_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4486_ (.A1(_0643_),
    .A2(_0649_),
    .B(_0642_),
    .ZN(_0924_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4487_ (.A1(_0614_),
    .A2(_0637_),
    .B1(_0639_),
    .B2(_0640_),
    .ZN(_0925_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4488_ (.A1(\r[14] ),
    .A2(net69),
    .ZN(_0926_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4489_ (.A1(\r[14] ),
    .A2(net78),
    .ZN(_0927_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4490_ (.A1(_0637_),
    .A2(_0927_),
    .Z(_0928_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4491_ (.A1(net148),
    .A2(\r[15] ),
    .ZN(_0929_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4492_ (.A1(_0637_),
    .A2(_0927_),
    .A3(_0929_),
    .ZN(_0930_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4493_ (.A1(_0925_),
    .A2(_0930_),
    .ZN(_0931_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4494_ (.A1(_0925_),
    .A2(_0930_),
    .ZN(_0932_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4495_ (.A1(\r[10] ),
    .A2(net51),
    .ZN(_0933_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4496_ (.A1(net107),
    .A2(net65),
    .ZN(_0934_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4497_ (.A1(net107),
    .A2(net67),
    .ZN(_0935_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4498_ (.A1(_0644_),
    .A2(_0935_),
    .Z(_0936_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4499_ (.A1(\r[10] ),
    .A2(net51),
    .A3(_0936_),
    .ZN(_0937_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4500_ (.A1(_0933_),
    .A2(_0936_),
    .ZN(_0938_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4501_ (.I(_0938_),
    .ZN(_0939_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4502_ (.A1(_0932_),
    .A2(_0938_),
    .ZN(_0940_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4503_ (.A1(_0924_),
    .A2(_0940_),
    .Z(_0941_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4504_ (.A1(_0924_),
    .A2(_0940_),
    .ZN(_0942_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4505_ (.A1(_0941_),
    .A2(_0942_),
    .ZN(_0943_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4506_ (.A1(_0923_),
    .A2(_0943_),
    .Z(_0944_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4507_ (.A1(_0918_),
    .A2(_0944_),
    .ZN(_0945_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4508_ (.A1(_0917_),
    .A2(_0944_),
    .Z(_0946_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4509_ (.A1(_0633_),
    .A2(_0946_),
    .Z(_0947_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4510_ (.A1(_0633_),
    .A2(_0946_),
    .ZN(_0948_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4511_ (.A1(_0947_),
    .A2(_0948_),
    .ZN(_0949_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4512_ (.A1(_0916_),
    .A2(_0949_),
    .ZN(_0950_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4513_ (.A1(_0916_),
    .A2(_0949_),
    .ZN(_0951_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4514_ (.A1(_0914_),
    .A2(_0916_),
    .A3(_0949_),
    .ZN(_0952_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _4515_ (.I0(_0897_),
    .I1(_0952_),
    .S(net57),
    .Z(_0953_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4516_ (.A1(net57),
    .A2(_0908_),
    .ZN(_0954_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _4517_ (.A1(_2768_),
    .A2(_0901_),
    .B(_0902_),
    .C(_0954_),
    .ZN(_0955_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4518_ (.A1(net56),
    .A2(_0910_),
    .ZN(_0956_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4519_ (.A1(_2862_),
    .A2(_0899_),
    .B(_0956_),
    .ZN(_0957_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4520_ (.A1(_0906_),
    .A2(_0957_),
    .ZN(_0958_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _4521_ (.A1(_2780_),
    .A2(_0953_),
    .B(_0955_),
    .C(_0958_),
    .ZN(\dot__t[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _4522_ (.A1(net4),
    .A2(_0951_),
    .B(_0950_),
    .ZN(_0959_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4523_ (.A1(_0923_),
    .A2(_0943_),
    .B(_0941_),
    .ZN(_0960_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4524_ (.I(_0960_),
    .ZN(_0961_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4525_ (.A1(_0644_),
    .A2(_0935_),
    .B(_0937_),
    .ZN(_0962_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4526_ (.A1(\r[9] ),
    .A2(_0590_),
    .B1(net49),
    .B2(\r[10] ),
    .ZN(_0963_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4527_ (.I(_0963_),
    .ZN(_0964_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4528_ (.A1(_0962_),
    .A2(_0964_),
    .ZN(_0965_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4529_ (.A1(_0962_),
    .A2(_0963_),
    .ZN(_0966_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4530_ (.A1(_0932_),
    .A2(_0939_),
    .B(_0931_),
    .ZN(_0967_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4531_ (.I(_0967_),
    .ZN(_0968_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4532_ (.A1(_0638_),
    .A2(_0926_),
    .B1(_0928_),
    .B2(_0929_),
    .ZN(_0969_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4533_ (.A1(\r[15] ),
    .A2(net69),
    .ZN(_0970_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4534_ (.A1(\r[15] ),
    .A2(net78),
    .ZN(_0971_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4535_ (.A1(_0926_),
    .A2(_0971_),
    .Z(_0972_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4536_ (.A1(net148),
    .A2(\r[16] ),
    .ZN(_0973_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4537_ (.A1(_0926_),
    .A2(_0971_),
    .A3(_0973_),
    .ZN(_0974_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4538_ (.A1(_0969_),
    .A2(_0974_),
    .ZN(_0975_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4539_ (.A1(_0969_),
    .A2(_0974_),
    .ZN(_0976_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4540_ (.A1(\r[13] ),
    .A2(net65),
    .ZN(_0977_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4541_ (.A1(\r[13] ),
    .A2(net67),
    .ZN(_0978_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4542_ (.A1(_0934_),
    .A2(_0978_),
    .Z(_0979_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4543_ (.A1(\r[11] ),
    .A2(net53),
    .ZN(_0980_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4544_ (.A1(_0934_),
    .A2(_0978_),
    .A3(_0980_),
    .ZN(_0981_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4545_ (.I(_0981_),
    .ZN(_0982_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4546_ (.A1(_0976_),
    .A2(_0982_),
    .ZN(_0983_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4547_ (.A1(_0968_),
    .A2(_0983_),
    .ZN(_0984_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4548_ (.A1(_0967_),
    .A2(_0983_),
    .Z(_0985_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4549_ (.I(_0985_),
    .ZN(_0986_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4550_ (.A1(_0966_),
    .A2(_0985_),
    .ZN(_0987_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4551_ (.A1(_0961_),
    .A2(_0987_),
    .ZN(_0988_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4552_ (.A1(_0960_),
    .A2(_0987_),
    .Z(_0989_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4553_ (.A1(_0922_),
    .A2(_0989_),
    .Z(_0990_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4554_ (.A1(_0922_),
    .A2(_0989_),
    .ZN(_0991_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4555_ (.A1(_0990_),
    .A2(_0991_),
    .ZN(_0992_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4556_ (.A1(_0945_),
    .A2(_0947_),
    .B(_0992_),
    .ZN(_0993_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4557_ (.I(_0993_),
    .ZN(_0994_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4558_ (.A1(_0945_),
    .A2(_0947_),
    .A3(_0992_),
    .ZN(_0995_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4559_ (.A1(_0994_),
    .A2(_0995_),
    .ZN(_0996_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4560_ (.A1(_0959_),
    .A2(_0996_),
    .ZN(_0997_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _4561_ (.I0(_0952_),
    .I1(_0997_),
    .S(net57),
    .Z(_0998_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4562_ (.A1(_0903_),
    .A2(_0911_),
    .Z(_0999_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai221_1 _4563_ (.A1(_0900_),
    .A2(_0907_),
    .B1(_0998_),
    .B2(_2780_),
    .C(_0999_),
    .ZN(\dot__t[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4564_ (.A1(_0966_),
    .A2(_0986_),
    .B(_0984_),
    .ZN(_1000_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4565_ (.I(_1000_),
    .ZN(_1001_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4566_ (.A1(_0935_),
    .A2(_0977_),
    .B1(_0979_),
    .B2(_0980_),
    .ZN(_1002_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4567_ (.A1(\r[10] ),
    .A2(net50),
    .B1(net48),
    .B2(\r[11] ),
    .ZN(_1003_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4568_ (.I(_1003_),
    .ZN(_1004_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4569_ (.A1(_1002_),
    .A2(_1004_),
    .ZN(_1005_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4570_ (.A1(_1002_),
    .A2(_1003_),
    .ZN(_1006_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4571_ (.A1(_0976_),
    .A2(_0982_),
    .B(_0975_),
    .ZN(_1007_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4572_ (.A1(_0927_),
    .A2(_0970_),
    .B1(_0972_),
    .B2(_0973_),
    .ZN(_1008_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4573_ (.A1(\r[16] ),
    .A2(net69),
    .ZN(_1009_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4574_ (.A1(\r[16] ),
    .A2(net78),
    .ZN(_1010_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4575_ (.A1(_0970_),
    .A2(_1010_),
    .Z(_1011_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4576_ (.A1(net148),
    .A2(\r[17] ),
    .ZN(_1012_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4577_ (.A1(_0970_),
    .A2(_1010_),
    .A3(_1012_),
    .ZN(_1013_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4578_ (.A1(_1008_),
    .A2(_1013_),
    .ZN(_1014_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4579_ (.A1(_1008_),
    .A2(_1013_),
    .ZN(_1015_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4580_ (.A1(net107),
    .A2(net53),
    .ZN(_1016_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4581_ (.A1(\r[14] ),
    .A2(net65),
    .ZN(_1017_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4582_ (.A1(\r[14] ),
    .A2(net67),
    .ZN(_1018_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4583_ (.A1(_0977_),
    .A2(_1018_),
    .Z(_1019_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4584_ (.A1(net107),
    .A2(net53),
    .A3(_1019_),
    .ZN(_1020_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4585_ (.A1(_1016_),
    .A2(_1019_),
    .ZN(_1021_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4586_ (.I(_1021_),
    .ZN(_1022_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4587_ (.A1(_1015_),
    .A2(_1021_),
    .ZN(_1023_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4588_ (.A1(_1007_),
    .A2(_1023_),
    .Z(_1024_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4589_ (.A1(_1007_),
    .A2(_1023_),
    .ZN(_1025_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4590_ (.A1(_1024_),
    .A2(_1025_),
    .ZN(_1026_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4591_ (.A1(_1006_),
    .A2(_1026_),
    .Z(_1027_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4592_ (.A1(_1001_),
    .A2(_1027_),
    .ZN(_1028_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4593_ (.A1(_1001_),
    .A2(_1027_),
    .ZN(_1029_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4594_ (.A1(_0965_),
    .A2(_1000_),
    .A3(_1027_),
    .ZN(_1030_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4595_ (.A1(_0988_),
    .A2(_0990_),
    .ZN(_1031_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4596_ (.A1(_0988_),
    .A2(_0990_),
    .B(_1030_),
    .ZN(_1032_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4597_ (.A1(_0988_),
    .A2(_0990_),
    .A3(_1030_),
    .ZN(_1033_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4598_ (.A1(_1030_),
    .A2(_1031_),
    .Z(_1034_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4599_ (.A1(_0959_),
    .A2(_0996_),
    .B(_0994_),
    .ZN(_1035_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4600_ (.A1(_1034_),
    .A2(_1035_),
    .ZN(_1036_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4601_ (.A1(net57),
    .A2(_0997_),
    .ZN(_1037_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4602_ (.A1(net57),
    .A2(_1036_),
    .B(_1037_),
    .ZN(_1038_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4603_ (.A1(_0902_),
    .A2(_0957_),
    .ZN(_1039_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai221_1 _4604_ (.A1(_0907_),
    .A2(_0953_),
    .B1(_1038_),
    .B2(_2780_),
    .C(_1039_),
    .ZN(\dot__t[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4605_ (.A1(_1006_),
    .A2(_1026_),
    .B(_1024_),
    .ZN(_1040_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4606_ (.I(_1040_),
    .ZN(_1041_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4607_ (.A1(_0977_),
    .A2(_1018_),
    .B(_1020_),
    .ZN(_1042_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4608_ (.A1(\r[11] ),
    .A2(net50),
    .B1(net49),
    .B2(\r[12] ),
    .ZN(_1043_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4609_ (.I(_1043_),
    .ZN(_1044_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4610_ (.A1(_1042_),
    .A2(_1044_),
    .ZN(_1045_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4611_ (.I(_1045_),
    .ZN(_1046_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4612_ (.A1(_1042_),
    .A2(_1043_),
    .ZN(_1047_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4613_ (.A1(_1015_),
    .A2(_1022_),
    .B(_1014_),
    .ZN(_1048_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4614_ (.I(_1048_),
    .ZN(_1049_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4615_ (.A1(_0971_),
    .A2(_1009_),
    .B1(_1011_),
    .B2(_1012_),
    .ZN(_1050_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4616_ (.A1(net148),
    .A2(\r[18] ),
    .ZN(_1051_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4617_ (.A1(\r[17] ),
    .A2(net69),
    .ZN(_1052_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4618_ (.A1(\r[17] ),
    .A2(net78),
    .ZN(_1053_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4619_ (.A1(_1009_),
    .A2(_1053_),
    .Z(_1054_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4620_ (.A1(_1009_),
    .A2(_1051_),
    .A3(_1053_),
    .ZN(_1055_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4621_ (.A1(_1050_),
    .A2(_1055_),
    .ZN(_1056_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4622_ (.A1(_1050_),
    .A2(_1055_),
    .ZN(_1057_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4623_ (.A1(\r[13] ),
    .A2(net53),
    .ZN(_1058_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4624_ (.A1(\r[15] ),
    .A2(net65),
    .ZN(_1059_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4625_ (.A1(\r[15] ),
    .A2(net67),
    .ZN(_1060_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4626_ (.A1(_1017_),
    .A2(_1060_),
    .Z(_1061_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4627_ (.A1(_1017_),
    .A2(_1058_),
    .A3(_1060_),
    .ZN(_1062_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4628_ (.I(_1062_),
    .ZN(_1063_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4629_ (.A1(_1057_),
    .A2(_1063_),
    .ZN(_1064_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4630_ (.A1(_1049_),
    .A2(_1064_),
    .ZN(_1065_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4631_ (.A1(_1048_),
    .A2(_1064_),
    .Z(_1066_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4632_ (.I(_1066_),
    .ZN(_1067_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4633_ (.A1(_1047_),
    .A2(_1066_),
    .ZN(_1068_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4634_ (.A1(_1041_),
    .A2(_1068_),
    .ZN(_1069_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4635_ (.A1(_1040_),
    .A2(_1068_),
    .Z(_1070_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4636_ (.A1(_1005_),
    .A2(_1070_),
    .Z(_1071_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4637_ (.A1(_0965_),
    .A2(_1029_),
    .B(_1028_),
    .ZN(_1072_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4638_ (.A1(_1071_),
    .A2(_1072_),
    .Z(_1073_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4639_ (.A1(_1071_),
    .A2(_1072_),
    .ZN(_1074_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4640_ (.I(_1074_),
    .ZN(_1075_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4641_ (.A1(_0993_),
    .A2(_1032_),
    .B(_1033_),
    .ZN(_1076_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _4642_ (.A1(_0959_),
    .A2(_0996_),
    .A3(_1034_),
    .B(_1076_),
    .ZN(_1077_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4643_ (.A1(_1074_),
    .A2(_1077_),
    .ZN(_1078_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _4644_ (.I0(_1036_),
    .I1(_1078_),
    .S(_2861_),
    .Z(_1079_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4645_ (.A1(_2780_),
    .A2(_1079_),
    .ZN(_1080_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _4646_ (.A1(_0900_),
    .A2(_0902_),
    .B1(_0906_),
    .B2(_0998_),
    .C(_1080_),
    .ZN(\dot__t[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4647_ (.A1(_2861_),
    .A2(_1078_),
    .Z(_1081_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4648_ (.A1(_1047_),
    .A2(_1067_),
    .B(_1065_),
    .ZN(_1082_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4649_ (.A1(_1057_),
    .A2(_1063_),
    .B(_1056_),
    .ZN(_1083_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4650_ (.A1(_1010_),
    .A2(_1052_),
    .B1(_1054_),
    .B2(_1051_),
    .ZN(_1084_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4651_ (.A1(net148),
    .A2(\r[19] ),
    .ZN(_1085_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4652_ (.A1(\r[18] ),
    .A2(net69),
    .ZN(_1086_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4653_ (.A1(\r[18] ),
    .A2(net79),
    .ZN(_1087_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4654_ (.A1(_1052_),
    .A2(_1087_),
    .Z(_1088_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4655_ (.A1(_1052_),
    .A2(_1085_),
    .A3(_1087_),
    .ZN(_1089_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4656_ (.A1(_1084_),
    .A2(_1089_),
    .ZN(_1090_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4657_ (.A1(_1084_),
    .A2(_1089_),
    .Z(_1091_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4658_ (.A1(\r[14] ),
    .A2(net51),
    .ZN(_1092_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4659_ (.A1(\r[16] ),
    .A2(net65),
    .ZN(_1093_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4660_ (.A1(\r[16] ),
    .A2(net67),
    .ZN(_1094_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4661_ (.A1(_1059_),
    .A2(_1094_),
    .Z(_1095_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4662_ (.A1(\r[14] ),
    .A2(net51),
    .A3(_1095_),
    .ZN(_1096_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4663_ (.A1(_1092_),
    .A2(_1095_),
    .ZN(_1097_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4664_ (.A1(_1091_),
    .A2(_1097_),
    .ZN(_1098_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4665_ (.A1(_1091_),
    .A2(_1097_),
    .ZN(_1099_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4666_ (.I(_1099_),
    .ZN(_1100_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4667_ (.A1(_1083_),
    .A2(_1100_),
    .ZN(_1101_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4668_ (.A1(_1083_),
    .A2(_1099_),
    .ZN(_1102_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4669_ (.A1(_1018_),
    .A2(_1059_),
    .B1(_1061_),
    .B2(_1058_),
    .ZN(_1103_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4670_ (.A1(\r[12] ),
    .A2(net50),
    .B1(net49),
    .B2(\r[13] ),
    .ZN(_1104_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4671_ (.I(_1104_),
    .ZN(_1105_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4672_ (.A1(_1103_),
    .A2(_1105_),
    .ZN(_1106_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4673_ (.A1(_1103_),
    .A2(_1104_),
    .ZN(_1107_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4674_ (.A1(_1102_),
    .A2(_1107_),
    .ZN(_1108_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4675_ (.A1(_1102_),
    .A2(_1107_),
    .ZN(_1109_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4676_ (.A1(_1082_),
    .A2(_1109_),
    .ZN(_1110_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4677_ (.A1(_1082_),
    .A2(_1109_),
    .ZN(_1111_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4678_ (.A1(_1045_),
    .A2(_1082_),
    .A3(_1109_),
    .ZN(_1112_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4679_ (.A1(_1005_),
    .A2(_1070_),
    .B(_1069_),
    .ZN(_1113_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4680_ (.A1(_1112_),
    .A2(_1113_),
    .ZN(_1114_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4681_ (.A1(_1112_),
    .A2(_1113_),
    .Z(_1115_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4682_ (.A1(_1114_),
    .A2(_1115_),
    .ZN(_1116_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4683_ (.A1(_1075_),
    .A2(_1077_),
    .B(_1073_),
    .ZN(_1117_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4684_ (.A1(_1116_),
    .A2(_1117_),
    .Z(_1118_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4685_ (.A1(_0902_),
    .A2(_0953_),
    .ZN(_1119_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _4686_ (.A1(net88),
    .A2(_2770_),
    .A3(_1078_),
    .B(_1119_),
    .ZN(_1120_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4687_ (.A1(_0906_),
    .A2(_1038_),
    .B(_1120_),
    .ZN(\dot__t[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4688_ (.A1(_0907_),
    .A2(_1079_),
    .B1(_1118_),
    .B2(_2780_),
    .ZN(_1121_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4689_ (.A1(_0902_),
    .A2(_0998_),
    .B(_1121_),
    .ZN(\dot__t[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _4690_ (.A1(_2862_),
    .A2(_1118_),
    .B(_1081_),
    .C(_0906_),
    .ZN(_1122_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4691_ (.A1(_1074_),
    .A2(_1116_),
    .ZN(_1123_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4692_ (.A1(_1073_),
    .A2(_1115_),
    .B1(_1123_),
    .B2(_1077_),
    .ZN(_1124_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4693_ (.A1(_1114_),
    .A2(_1124_),
    .ZN(_1125_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4694_ (.A1(net141),
    .A2(\r[19] ),
    .ZN(_1126_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4695_ (.A1(_1053_),
    .A2(_1086_),
    .B1(_1088_),
    .B2(_1085_),
    .ZN(_1127_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4696_ (.A1(\r[17] ),
    .A2(net67),
    .ZN(_1128_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _4697_ (.A1(_1093_),
    .A2(_1127_),
    .A3(_1128_),
    .Z(_1129_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4698_ (.A1(_1086_),
    .A2(_1126_),
    .A3(_1129_),
    .ZN(_1130_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4699_ (.A1(\r[15] ),
    .A2(net51),
    .ZN(_1131_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4700_ (.A1(\r[13] ),
    .A2(_0590_),
    .B1(net49),
    .B2(\r[14] ),
    .ZN(_1132_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4701_ (.A1(_1130_),
    .A2(_1131_),
    .A3(_1132_),
    .ZN(_1133_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4702_ (.A1(_1090_),
    .A2(_1098_),
    .ZN(_1134_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4703_ (.A1(_1059_),
    .A2(_1094_),
    .B(_1096_),
    .ZN(_1135_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4704_ (.A1(_1133_),
    .A2(_1134_),
    .A3(_1135_),
    .ZN(_1136_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4705_ (.A1(_1101_),
    .A2(_1108_),
    .ZN(_1137_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4706_ (.A1(_1106_),
    .A2(_1137_),
    .Z(_1138_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4707_ (.A1(_1136_),
    .A2(_1138_),
    .ZN(_1139_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4708_ (.A1(_1046_),
    .A2(_1111_),
    .B(_1110_),
    .ZN(_1140_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4709_ (.A1(_1125_),
    .A2(_1139_),
    .A3(_1140_),
    .ZN(_1141_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai221_1 _4710_ (.A1(_0903_),
    .A2(_1038_),
    .B1(_1141_),
    .B2(_2780_),
    .C(_1122_),
    .ZN(\dot__t[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4711_ (.A1(net114),
    .A2(\pp_x_sq[7] ),
    .ZN(_1142_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4712_ (.A1(net138),
    .A2(\pp_x_sq[10] ),
    .ZN(_1143_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4713_ (.A1(net145),
    .A2(\pp_x_sq[9] ),
    .ZN(_1144_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4714_ (.A1(net145),
    .A2(\pp_x_sq[10] ),
    .ZN(_1145_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4715_ (.A1(net138),
    .A2(\pp_x_sq[9] ),
    .ZN(_1146_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4716_ (.A1(net133),
    .A2(\pp_x_sq[8] ),
    .ZN(_1147_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4717_ (.A1(net145),
    .A2(\pp_x_sq[10] ),
    .B1(\pp_x_sq[9] ),
    .B2(net138),
    .ZN(_1148_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4718_ (.A1(_1143_),
    .A2(_1144_),
    .B1(_1147_),
    .B2(_1148_),
    .ZN(_1149_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4719_ (.A1(net133),
    .A2(\pp_x_sq[9] ),
    .ZN(_1150_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4720_ (.A1(net138),
    .A2(\pp_x_sq[11] ),
    .ZN(_1151_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4721_ (.A1(net145),
    .A2(\pp_x_sq[11] ),
    .ZN(_1152_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4722_ (.A1(net145),
    .A2(\pp_x_sq[11] ),
    .B1(\pp_x_sq[10] ),
    .B2(net138),
    .ZN(_1153_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4723_ (.A1(_1143_),
    .A2(_1150_),
    .A3(_1152_),
    .ZN(_1154_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4724_ (.A1(_1149_),
    .A2(_1154_),
    .ZN(_1155_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4725_ (.A1(net119),
    .A2(\pp_x_sq[6] ),
    .ZN(_1156_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4726_ (.A1(net124),
    .A2(\pp_x_sq[8] ),
    .ZN(_1157_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4727_ (.A1(net128),
    .A2(\pp_x_sq[7] ),
    .ZN(_1158_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4728_ (.A1(net128),
    .A2(\pp_x_sq[8] ),
    .ZN(_1159_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4729_ (.A1(net124),
    .A2(\pp_x_sq[7] ),
    .ZN(_1160_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4730_ (.A1(_1159_),
    .A2(_1160_),
    .ZN(_1161_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4731_ (.A1(_1156_),
    .A2(_1161_),
    .ZN(_1162_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4732_ (.A1(_1149_),
    .A2(_1154_),
    .ZN(_1163_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4733_ (.A1(_1162_),
    .A2(_1163_),
    .B(_1155_),
    .ZN(_1164_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4734_ (.A1(net124),
    .A2(\pp_x_sq[9] ),
    .ZN(_1165_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4735_ (.A1(net128),
    .A2(\pp_x_sq[9] ),
    .ZN(_1166_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4736_ (.A1(_1157_),
    .A2(_1166_),
    .Z(_1167_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4737_ (.A1(net119),
    .A2(\pp_x_sq[7] ),
    .ZN(_1168_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4738_ (.A1(_1157_),
    .A2(_1166_),
    .A3(_1168_),
    .ZN(_1169_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4739_ (.A1(_1145_),
    .A2(_1151_),
    .B1(_1153_),
    .B2(_1150_),
    .ZN(_1170_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4740_ (.A1(net133),
    .A2(\pp_x_sq[10] ),
    .ZN(_1171_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4741_ (.A1(net138),
    .A2(\pp_x_sq[12] ),
    .ZN(_1172_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4742_ (.A1(net146),
    .A2(\pp_x_sq[12] ),
    .ZN(_1173_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4743_ (.A1(_1151_),
    .A2(_1173_),
    .Z(_1174_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4744_ (.A1(_1151_),
    .A2(_1171_),
    .A3(_1173_),
    .ZN(_1175_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4745_ (.A1(_1170_),
    .A2(_1175_),
    .ZN(_1176_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4746_ (.A1(_1170_),
    .A2(_1175_),
    .Z(_1177_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4747_ (.A1(_1169_),
    .A2(_1177_),
    .ZN(_1178_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4748_ (.A1(_1169_),
    .A2(_1177_),
    .ZN(_1179_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4749_ (.I(_1179_),
    .ZN(_1180_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4750_ (.A1(_1164_),
    .A2(_1180_),
    .ZN(_1181_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4751_ (.A1(_1157_),
    .A2(_1158_),
    .B1(_1161_),
    .B2(_1156_),
    .ZN(_1182_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4752_ (.I(_1182_),
    .ZN(_1183_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4753_ (.A1(_1164_),
    .A2(_1179_),
    .Z(_1184_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4754_ (.A1(_1183_),
    .A2(_1184_),
    .B(_1181_),
    .ZN(_1185_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4755_ (.A1(_1159_),
    .A2(_1165_),
    .B1(_1167_),
    .B2(_1168_),
    .ZN(_1186_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4756_ (.I(_1186_),
    .ZN(_1187_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4757_ (.A1(_1176_),
    .A2(_1178_),
    .ZN(_1188_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4758_ (.A1(net119),
    .A2(\pp_x_sq[8] ),
    .ZN(_1189_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4759_ (.A1(net125),
    .A2(\pp_x_sq[10] ),
    .ZN(_1190_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4760_ (.A1(net128),
    .A2(\pp_x_sq[10] ),
    .ZN(_1191_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4761_ (.A1(_1165_),
    .A2(_1191_),
    .ZN(_1192_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4762_ (.A1(_1189_),
    .A2(_1192_),
    .Z(_1193_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4763_ (.A1(_1152_),
    .A2(_1172_),
    .B1(_1174_),
    .B2(_1171_),
    .ZN(_1194_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4764_ (.A1(net132),
    .A2(\pp_x_sq[11] ),
    .ZN(_1195_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4765_ (.A1(net140),
    .A2(\pp_x_sq[13] ),
    .ZN(_1196_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4766_ (.A1(net145),
    .A2(\pp_x_sq[13] ),
    .ZN(_1197_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4767_ (.A1(_1172_),
    .A2(_1197_),
    .Z(_1198_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4768_ (.A1(net132),
    .A2(\pp_x_sq[11] ),
    .A3(_1198_),
    .ZN(_1199_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4769_ (.A1(_1195_),
    .A2(_1198_),
    .ZN(_1200_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4770_ (.A1(_1194_),
    .A2(_1200_),
    .ZN(_1201_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4771_ (.A1(_1194_),
    .A2(_1200_),
    .Z(_1202_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4772_ (.A1(_1193_),
    .A2(_1201_),
    .A3(_1202_),
    .ZN(_1203_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4773_ (.A1(_1193_),
    .A2(_1194_),
    .A3(_1200_),
    .ZN(_1204_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4774_ (.I(_1204_),
    .ZN(_1205_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4775_ (.A1(_1188_),
    .A2(_1205_),
    .ZN(_1206_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4776_ (.A1(_1188_),
    .A2(_1205_),
    .ZN(_1207_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4777_ (.A1(_1186_),
    .A2(_1207_),
    .ZN(_1208_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4778_ (.A1(_1185_),
    .A2(_1208_),
    .ZN(_1209_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4779_ (.A1(_1185_),
    .A2(_1208_),
    .Z(_1210_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4780_ (.A1(net114),
    .A2(\pp_x_sq[7] ),
    .A3(_1210_),
    .ZN(_1211_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4781_ (.A1(_1142_),
    .A2(_1210_),
    .ZN(_1212_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4782_ (.A1(net145),
    .A2(\pp_x_sq[8] ),
    .ZN(_1213_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4783_ (.A1(net138),
    .A2(\pp_x_sq[8] ),
    .ZN(_1214_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4784_ (.A1(net133),
    .A2(\pp_x_sq[7] ),
    .ZN(_1215_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4785_ (.A1(net145),
    .A2(\pp_x_sq[9] ),
    .B1(\pp_x_sq[8] ),
    .B2(net138),
    .ZN(_1216_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4786_ (.A1(_1146_),
    .A2(_1213_),
    .B1(_1215_),
    .B2(_1216_),
    .ZN(_1217_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4787_ (.A1(_1145_),
    .A2(_1146_),
    .A3(_1147_),
    .ZN(_1218_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4788_ (.A1(_1217_),
    .A2(_1218_),
    .ZN(_1219_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4789_ (.A1(net119),
    .A2(\pp_x_sq[5] ),
    .ZN(_1220_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4790_ (.A1(net128),
    .A2(\pp_x_sq[6] ),
    .ZN(_1221_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4791_ (.A1(net124),
    .A2(\pp_x_sq[6] ),
    .ZN(_1222_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4792_ (.A1(_1160_),
    .A2(_1221_),
    .ZN(_1223_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4793_ (.A1(_1158_),
    .A2(_1222_),
    .ZN(_1224_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4794_ (.A1(_1220_),
    .A2(_1224_),
    .ZN(_1225_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4795_ (.A1(_1220_),
    .A2(_1224_),
    .ZN(_1226_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4796_ (.A1(_1217_),
    .A2(_1218_),
    .ZN(_1227_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4797_ (.A1(_1226_),
    .A2(_1227_),
    .B(_1219_),
    .ZN(_1228_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4798_ (.A1(_1162_),
    .A2(_1163_),
    .Z(_1229_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4799_ (.A1(_1228_),
    .A2(_1229_),
    .ZN(_1230_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4800_ (.A1(_1223_),
    .A2(_1225_),
    .ZN(_1231_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4801_ (.A1(_1228_),
    .A2(_1229_),
    .ZN(_1232_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4802_ (.A1(_1231_),
    .A2(_1232_),
    .B(_1230_),
    .ZN(_1233_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4803_ (.A1(_1182_),
    .A2(_1184_),
    .ZN(_1234_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4804_ (.A1(_1233_),
    .A2(_1234_),
    .ZN(_1235_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4805_ (.A1(net114),
    .A2(\pp_x_sq[6] ),
    .ZN(_1236_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4806_ (.A1(_1233_),
    .A2(_1234_),
    .ZN(_1237_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4807_ (.A1(_1236_),
    .A2(_1237_),
    .B(_1235_),
    .ZN(_1238_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4808_ (.A1(_1212_),
    .A2(_1238_),
    .ZN(_1239_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4809_ (.I(_1239_),
    .ZN(_1240_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4810_ (.A1(_1212_),
    .A2(_1238_),
    .ZN(_1241_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4811_ (.A1(net145),
    .A2(\pp_x_sq[7] ),
    .ZN(_1242_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4812_ (.A1(net138),
    .A2(\pp_x_sq[7] ),
    .ZN(_1243_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4813_ (.A1(net133),
    .A2(\pp_x_sq[6] ),
    .ZN(_1244_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4814_ (.A1(net145),
    .A2(\pp_x_sq[8] ),
    .B1(\pp_x_sq[7] ),
    .B2(net138),
    .ZN(_1245_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4815_ (.A1(_1214_),
    .A2(_1242_),
    .B1(_1244_),
    .B2(_1245_),
    .ZN(_1246_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4816_ (.A1(_1144_),
    .A2(_1214_),
    .A3(_1215_),
    .ZN(_1247_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4817_ (.A1(_1246_),
    .A2(_1247_),
    .ZN(_1248_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4818_ (.A1(net119),
    .A2(\pp_x_sq[4] ),
    .ZN(_1249_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4819_ (.A1(net128),
    .A2(\pp_x_sq[5] ),
    .ZN(_1250_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4820_ (.A1(net124),
    .A2(\pp_x_sq[5] ),
    .ZN(_1251_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4821_ (.A1(_1221_),
    .A2(_1251_),
    .Z(_1252_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4822_ (.A1(net119),
    .A2(\pp_x_sq[4] ),
    .A3(_1252_),
    .ZN(_1253_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4823_ (.A1(_1249_),
    .A2(_1252_),
    .Z(_1254_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4824_ (.A1(_1246_),
    .A2(_1247_),
    .ZN(_1255_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4825_ (.A1(_1254_),
    .A2(_1255_),
    .B(_1248_),
    .ZN(_1256_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4826_ (.A1(_1226_),
    .A2(_1227_),
    .Z(_1257_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4827_ (.A1(_1256_),
    .A2(_1257_),
    .ZN(_1258_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4828_ (.A1(_1221_),
    .A2(_1251_),
    .B(_1253_),
    .ZN(_1259_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4829_ (.I(_1259_),
    .ZN(_1260_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4830_ (.A1(_1256_),
    .A2(_1257_),
    .ZN(_1261_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4831_ (.A1(_1260_),
    .A2(_1261_),
    .B(_1258_),
    .ZN(_1262_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4832_ (.A1(_1231_),
    .A2(_1232_),
    .Z(_1263_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4833_ (.A1(_1262_),
    .A2(_1263_),
    .ZN(_1264_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4834_ (.A1(net114),
    .A2(\pp_x_sq[5] ),
    .ZN(_1265_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4835_ (.A1(_1262_),
    .A2(_1263_),
    .ZN(_1266_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4836_ (.A1(_1265_),
    .A2(_1266_),
    .B(_1264_),
    .ZN(_1267_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4837_ (.A1(_1236_),
    .A2(_1237_),
    .Z(_1268_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4838_ (.A1(_1267_),
    .A2(_1268_),
    .ZN(_1269_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4839_ (.A1(net114),
    .A2(\pp_x_sq[4] ),
    .ZN(_1270_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4840_ (.I(_1270_),
    .ZN(_1271_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4841_ (.A1(net146),
    .A2(\pp_x_sq[6] ),
    .ZN(_1272_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4842_ (.A1(net139),
    .A2(\pp_x_sq[6] ),
    .ZN(_1273_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4843_ (.A1(net133),
    .A2(\pp_x_sq[5] ),
    .ZN(_1274_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4844_ (.A1(net146),
    .A2(\pp_x_sq[7] ),
    .B1(\pp_x_sq[6] ),
    .B2(net139),
    .ZN(_1275_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4845_ (.A1(_1243_),
    .A2(_1272_),
    .B1(_1274_),
    .B2(_1275_),
    .ZN(_1276_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4846_ (.A1(_1213_),
    .A2(_1243_),
    .A3(_1244_),
    .ZN(_1277_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4847_ (.A1(_1276_),
    .A2(_1277_),
    .ZN(_1278_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4848_ (.A1(net129),
    .A2(\pp_x_sq[4] ),
    .ZN(_1279_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4849_ (.A1(net125),
    .A2(\pp_x_sq[4] ),
    .ZN(_1280_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4850_ (.A1(_1250_),
    .A2(_1280_),
    .Z(_1281_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4851_ (.A1(net119),
    .A2(\pp_x_sq[3] ),
    .ZN(_1282_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _4852_ (.A1(_1250_),
    .A2(_1280_),
    .A3(_1282_),
    .Z(_1283_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4853_ (.A1(_1276_),
    .A2(_1277_),
    .ZN(_1284_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4854_ (.A1(_1283_),
    .A2(_1284_),
    .B(_1278_),
    .ZN(_1285_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4855_ (.A1(_1254_),
    .A2(_1255_),
    .Z(_1286_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4856_ (.A1(_1285_),
    .A2(_1286_),
    .ZN(_1287_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4857_ (.A1(_1251_),
    .A2(_1279_),
    .B1(_1281_),
    .B2(_1282_),
    .ZN(_1288_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4858_ (.I(_1288_),
    .ZN(_1289_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4859_ (.A1(_1285_),
    .A2(_1286_),
    .ZN(_1290_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4860_ (.A1(_1289_),
    .A2(_1290_),
    .B(_1287_),
    .ZN(_1291_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4861_ (.A1(_1259_),
    .A2(_1261_),
    .ZN(_1292_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4862_ (.A1(_1291_),
    .A2(_1292_),
    .Z(_1293_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4863_ (.A1(_1291_),
    .A2(_1292_),
    .Z(_1294_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4864_ (.A1(_1271_),
    .A2(_1291_),
    .A3(_1292_),
    .ZN(_1295_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4865_ (.A1(net146),
    .A2(\pp_x_sq[5] ),
    .ZN(_1296_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4866_ (.A1(net139),
    .A2(\pp_x_sq[5] ),
    .ZN(_1297_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4867_ (.A1(net132),
    .A2(\pp_x_sq[4] ),
    .ZN(_1298_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4868_ (.A1(net146),
    .A2(\pp_x_sq[6] ),
    .B1(\pp_x_sq[5] ),
    .B2(net139),
    .ZN(_1299_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4869_ (.A1(_1273_),
    .A2(_1296_),
    .B1(_1298_),
    .B2(_1299_),
    .ZN(_1300_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4870_ (.A1(_1242_),
    .A2(_1273_),
    .A3(_1274_),
    .ZN(_1301_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4871_ (.A1(_1300_),
    .A2(_1301_),
    .ZN(_1302_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4872_ (.A1(net124),
    .A2(\pp_x_sq[3] ),
    .ZN(_1303_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4873_ (.A1(_1279_),
    .A2(_1303_),
    .Z(_1304_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4874_ (.A1(net120),
    .A2(\pp_x_sq[2] ),
    .ZN(_1305_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4875_ (.A1(net119),
    .A2(\pp_x_sq[2] ),
    .A3(_1304_),
    .ZN(_1306_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4876_ (.A1(_1304_),
    .A2(_1305_),
    .Z(_1307_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4877_ (.A1(_1300_),
    .A2(_1301_),
    .ZN(_1308_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4878_ (.A1(_1307_),
    .A2(_1308_),
    .B(_1302_),
    .ZN(_1309_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4879_ (.A1(_1283_),
    .A2(_1284_),
    .Z(_1310_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4880_ (.A1(_1309_),
    .A2(_1310_),
    .Z(_1311_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4881_ (.A1(_1279_),
    .A2(_1303_),
    .B(_1306_),
    .ZN(_1312_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4882_ (.A1(_1309_),
    .A2(_1310_),
    .Z(_1313_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4883_ (.A1(_1312_),
    .A2(_1313_),
    .B(_1311_),
    .ZN(_1314_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4884_ (.A1(_1289_),
    .A2(_1290_),
    .ZN(_1315_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4885_ (.A1(_1314_),
    .A2(_1315_),
    .ZN(_1316_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4886_ (.A1(net114),
    .A2(\pp_x_sq[3] ),
    .Z(_1317_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4887_ (.A1(_1314_),
    .A2(_1315_),
    .ZN(_1318_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4888_ (.A1(_1317_),
    .A2(_1318_),
    .B(_1316_),
    .ZN(_1319_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4889_ (.A1(_1295_),
    .A2(_1319_),
    .ZN(_1320_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4890_ (.A1(net114),
    .A2(\pp_x_sq[2] ),
    .Z(_1321_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4891_ (.A1(_1312_),
    .A2(_1313_),
    .ZN(_1322_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4892_ (.A1(net146),
    .A2(\pp_x_sq[4] ),
    .ZN(_1323_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4893_ (.A1(net139),
    .A2(\pp_x_sq[4] ),
    .ZN(_1324_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4894_ (.A1(net132),
    .A2(\pp_x_sq[3] ),
    .ZN(_1325_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4895_ (.A1(net146),
    .A2(\pp_x_sq[5] ),
    .B1(\pp_x_sq[4] ),
    .B2(net139),
    .ZN(_1326_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4896_ (.A1(_1297_),
    .A2(_1323_),
    .B1(_1325_),
    .B2(_1326_),
    .ZN(_1327_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4897_ (.A1(_1272_),
    .A2(_1297_),
    .A3(_1298_),
    .ZN(_1328_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4898_ (.A1(net128),
    .A2(\pp_x_sq[3] ),
    .B1(\pp_x_sq[2] ),
    .B2(net124),
    .ZN(_1329_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4899_ (.A1(net128),
    .A2(\pp_x_sq[2] ),
    .ZN(_1330_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4900_ (.A1(_1303_),
    .A2(_1330_),
    .ZN(_1331_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4901_ (.A1(_1329_),
    .A2(_1331_),
    .ZN(_1332_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4902_ (.A1(_1327_),
    .A2(_1328_),
    .Z(_1333_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4903_ (.A1(_1327_),
    .A2(_1328_),
    .B1(_1332_),
    .B2(_1333_),
    .ZN(_1334_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4904_ (.A1(_1307_),
    .A2(_1308_),
    .ZN(_1335_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4905_ (.A1(_1334_),
    .A2(_1335_),
    .ZN(_1336_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4906_ (.A1(_1334_),
    .A2(_1335_),
    .Z(_1337_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4907_ (.A1(_1331_),
    .A2(_1337_),
    .B(_1336_),
    .ZN(_1338_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4908_ (.A1(_1322_),
    .A2(_1338_),
    .ZN(_1339_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4909_ (.A1(_1322_),
    .A2(_1338_),
    .ZN(_1340_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4910_ (.A1(_1322_),
    .A2(_1338_),
    .Z(_1341_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4911_ (.A1(_1331_),
    .A2(_1337_),
    .ZN(_1342_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4912_ (.A1(net146),
    .A2(\pp_x_sq[3] ),
    .ZN(_1343_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4913_ (.A1(net141),
    .A2(\pp_x_sq[3] ),
    .ZN(_1344_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4914_ (.A1(net134),
    .A2(\pp_x_sq[2] ),
    .ZN(_1345_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4915_ (.A1(net146),
    .A2(\pp_x_sq[4] ),
    .B1(\pp_x_sq[3] ),
    .B2(net139),
    .ZN(_1346_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4916_ (.A1(_1324_),
    .A2(_1343_),
    .B1(_1345_),
    .B2(_1346_),
    .ZN(_1347_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4917_ (.A1(_1296_),
    .A2(_1324_),
    .A3(_1325_),
    .ZN(_1348_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4918_ (.A1(_1347_),
    .A2(_1348_),
    .ZN(_1349_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4919_ (.A1(net119),
    .A2(\pp_x_sq[0] ),
    .ZN(_1350_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4920_ (.A1(_1330_),
    .A2(_1350_),
    .ZN(_1351_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4921_ (.A1(net128),
    .A2(\pp_x_sq[2] ),
    .B1(\pp_x_sq[0] ),
    .B2(net120),
    .ZN(_1352_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4922_ (.A1(_1351_),
    .A2(_1352_),
    .ZN(_1353_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4923_ (.A1(_1347_),
    .A2(_1348_),
    .ZN(_1354_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _4924_ (.A1(_1351_),
    .A2(_1352_),
    .A3(_1354_),
    .B(_1349_),
    .ZN(_1355_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4925_ (.A1(_1332_),
    .A2(_1333_),
    .Z(_1356_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4926_ (.A1(_1355_),
    .A2(_1356_),
    .Z(_1357_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4927_ (.A1(_1355_),
    .A2(_1356_),
    .Z(_1358_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4928_ (.A1(_1351_),
    .A2(_1358_),
    .B(_1357_),
    .ZN(_1359_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4929_ (.A1(_1342_),
    .A2(_1359_),
    .ZN(_1360_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4930_ (.A1(net115),
    .A2(\pp_x_sq[0] ),
    .Z(_1361_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _4931_ (.A1(_1351_),
    .A2(_1355_),
    .A3(_1356_),
    .Z(_1362_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and4_1 _4932_ (.A1(net141),
    .A2(net150),
    .A3(\pp_x_sq[3] ),
    .A4(\pp_x_sq[2] ),
    .Z(_1363_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4933_ (.A1(_1323_),
    .A2(_1344_),
    .A3(_1345_),
    .ZN(_1364_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4934_ (.A1(_1363_),
    .A2(_1364_),
    .ZN(_1365_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _4935_ (.A1(net150),
    .A2(\pp_x_sq[3] ),
    .B1(\pp_x_sq[2] ),
    .B2(net141),
    .ZN(_1366_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai32_1 _4936_ (.A1(_2549_),
    .A2(_2552_),
    .A3(_1345_),
    .B1(_1363_),
    .B2(_1366_),
    .ZN(_1367_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4937_ (.A1(_2552_),
    .A2(_1345_),
    .B(_2549_),
    .ZN(_1368_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _4938_ (.A1(\pp_x_sq[0] ),
    .A2(_1367_),
    .A3(_1368_),
    .Z(_1369_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4939_ (.A1(net125),
    .A2(\pp_x_sq[0] ),
    .B(_1369_),
    .ZN(_1370_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4940_ (.A1(_1363_),
    .A2(_1364_),
    .ZN(_1371_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4941_ (.A1(net125),
    .A2(_1369_),
    .ZN(_1372_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _4942_ (.A1(_1365_),
    .A2(_1370_),
    .B(_1371_),
    .C(_1372_),
    .ZN(_1373_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4943_ (.A1(_1353_),
    .A2(_1354_),
    .ZN(_1374_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4944_ (.A1(_1371_),
    .A2(_1372_),
    .ZN(_1375_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _4945_ (.A1(_1361_),
    .A2(_1362_),
    .B1(_1373_),
    .B2(_1374_),
    .C(_1375_),
    .ZN(_1376_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4946_ (.A1(_1361_),
    .A2(_1362_),
    .ZN(_1377_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _4947_ (.A1(_1342_),
    .A2(_1359_),
    .B(_1376_),
    .C(_1377_),
    .ZN(_1378_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4948_ (.A1(_1321_),
    .A2(_1341_),
    .B1(_1360_),
    .B2(_1378_),
    .ZN(_1379_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _4949_ (.A1(_1314_),
    .A2(_1315_),
    .A3(_1317_),
    .Z(_1380_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _4950_ (.A1(_1321_),
    .A2(_1339_),
    .B(_1340_),
    .C(_1380_),
    .ZN(_1381_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4951_ (.A1(_1339_),
    .A2(_1380_),
    .ZN(_1382_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4952_ (.A1(_1271_),
    .A2(_1294_),
    .B(_1293_),
    .ZN(_1383_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4953_ (.A1(_1265_),
    .A2(_1266_),
    .ZN(_1384_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4954_ (.A1(_1383_),
    .A2(_1384_),
    .ZN(_1385_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _4955_ (.A1(_1295_),
    .A2(_1319_),
    .B1(_1379_),
    .B2(_1381_),
    .C(_1382_),
    .ZN(_1386_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4956_ (.A1(_1320_),
    .A2(_1386_),
    .B(_1385_),
    .ZN(_1387_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _4957_ (.A1(_1383_),
    .A2(_1384_),
    .ZN(_1388_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4958_ (.A1(_1267_),
    .A2(_1268_),
    .B(_1388_),
    .ZN(_1389_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _4959_ (.A1(_1387_),
    .A2(_1389_),
    .B(_1269_),
    .ZN(_1390_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _4960_ (.A1(_2543_),
    .A2(_0224_),
    .A3(net80),
    .ZN(_1391_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _4961_ (.A1(net111),
    .A2(_0225_),
    .A3(net71),
    .ZN(_1392_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _4962_ (.A1(_1387_),
    .A2(_1389_),
    .B(_1241_),
    .C(_1269_),
    .ZN(_1393_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4963_ (.A1(net114),
    .A2(\pp_x_sq[8] ),
    .ZN(_1394_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4964_ (.A1(_1187_),
    .A2(_1207_),
    .B(_1206_),
    .ZN(_1395_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _4965_ (.A1(_1166_),
    .A2(_1190_),
    .B1(_1192_),
    .B2(_1189_),
    .ZN(_1396_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4966_ (.I(_1396_),
    .ZN(_1397_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4967_ (.A1(_1201_),
    .A2(_1203_),
    .ZN(_1398_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4968_ (.A1(net119),
    .A2(\pp_x_sq[9] ),
    .ZN(_1399_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4969_ (.A1(net124),
    .A2(\pp_x_sq[11] ),
    .ZN(_1400_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4970_ (.A1(net128),
    .A2(\pp_x_sq[11] ),
    .ZN(_1401_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4971_ (.A1(_1190_),
    .A2(_1401_),
    .ZN(_1402_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4972_ (.A1(_1399_),
    .A2(_1402_),
    .Z(_1403_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4973_ (.A1(_1172_),
    .A2(_1197_),
    .B(_1199_),
    .ZN(_1404_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4974_ (.A1(net132),
    .A2(\pp_x_sq[12] ),
    .ZN(_1405_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4975_ (.A1(net140),
    .A2(\pp_x_sq[14] ),
    .ZN(_1406_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4976_ (.A1(net147),
    .A2(\pp_x_sq[14] ),
    .ZN(_1407_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _4977_ (.A1(_1196_),
    .A2(_1407_),
    .Z(_1408_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4978_ (.A1(_1196_),
    .A2(_1405_),
    .A3(_1407_),
    .ZN(_1409_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4979_ (.A1(_1404_),
    .A2(_1409_),
    .ZN(_1410_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _4980_ (.A1(_1404_),
    .A2(_1409_),
    .Z(_1411_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4981_ (.A1(_1403_),
    .A2(_1410_),
    .A3(_1411_),
    .ZN(_1412_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _4982_ (.A1(_1403_),
    .A2(_1404_),
    .A3(_1409_),
    .ZN(_1413_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4983_ (.I(_1413_),
    .ZN(_1414_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4984_ (.A1(_1398_),
    .A2(_1414_),
    .ZN(_1415_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4985_ (.A1(_1398_),
    .A2(_1414_),
    .ZN(_1416_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4986_ (.A1(_1396_),
    .A2(_1416_),
    .ZN(_1417_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4987_ (.A1(_1395_),
    .A2(_1417_),
    .ZN(_1418_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4988_ (.A1(_1395_),
    .A2(_1417_),
    .Z(_1419_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _4989_ (.A1(net114),
    .A2(\pp_x_sq[8] ),
    .A3(_1419_),
    .ZN(_1420_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _4990_ (.A1(_1394_),
    .A2(_1419_),
    .Z(_1421_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _4991_ (.I(_1421_),
    .ZN(_1422_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4992_ (.A1(_1209_),
    .A2(_1211_),
    .ZN(_1423_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4993_ (.A1(_1422_),
    .A2(_1423_),
    .ZN(_1424_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _4994_ (.A1(_1421_),
    .A2(_1423_),
    .ZN(_1425_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4995_ (.A1(_1240_),
    .A2(_1393_),
    .B(_1425_),
    .ZN(_1426_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4996_ (.A1(_1424_),
    .A2(_1426_),
    .ZN(_1427_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4997_ (.A1(_1418_),
    .A2(_1420_),
    .ZN(_1428_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _4998_ (.A1(net115),
    .A2(\pp_x_sq[9] ),
    .ZN(_1429_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _4999_ (.A1(_1397_),
    .A2(_1416_),
    .B(_1415_),
    .ZN(_1430_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5000_ (.A1(_1191_),
    .A2(_1400_),
    .B1(_1402_),
    .B2(_1399_),
    .ZN(_1431_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5001_ (.I(_1431_),
    .ZN(_1432_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5002_ (.A1(_1410_),
    .A2(_1412_),
    .ZN(_1433_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5003_ (.A1(_1197_),
    .A2(_1406_),
    .B1(_1408_),
    .B2(_1405_),
    .ZN(_1434_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5004_ (.A1(net147),
    .A2(\pp_x_sq[15] ),
    .ZN(_1435_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5005_ (.A1(net140),
    .A2(\pp_x_sq[15] ),
    .ZN(_1436_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5006_ (.A1(_1406_),
    .A2(_1435_),
    .Z(_1437_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5007_ (.A1(net132),
    .A2(\pp_x_sq[13] ),
    .ZN(_1438_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5008_ (.A1(net132),
    .A2(\pp_x_sq[13] ),
    .A3(_1437_),
    .ZN(_1439_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5009_ (.A1(_1437_),
    .A2(_1438_),
    .ZN(_1440_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5010_ (.A1(_1434_),
    .A2(_1440_),
    .ZN(_1441_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5011_ (.A1(_1434_),
    .A2(_1440_),
    .ZN(_1442_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5012_ (.I(_1442_),
    .ZN(_1443_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5013_ (.A1(net120),
    .A2(\pp_x_sq[10] ),
    .ZN(_1444_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5014_ (.A1(net124),
    .A2(\pp_x_sq[12] ),
    .ZN(_1445_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5015_ (.A1(net129),
    .A2(\pp_x_sq[12] ),
    .ZN(_1446_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5016_ (.A1(_1400_),
    .A2(_1446_),
    .ZN(_1447_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5017_ (.A1(_1444_),
    .A2(_1447_),
    .Z(_1448_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5018_ (.A1(_1443_),
    .A2(_1448_),
    .ZN(_1449_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5019_ (.A1(_1442_),
    .A2(_1448_),
    .Z(_1450_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5020_ (.I(_1450_),
    .ZN(_1451_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5021_ (.A1(_1433_),
    .A2(_1451_),
    .ZN(_1452_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5022_ (.A1(_1433_),
    .A2(_1451_),
    .ZN(_1453_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5023_ (.A1(_1431_),
    .A2(_1453_),
    .ZN(_1454_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5024_ (.A1(_1430_),
    .A2(_1454_),
    .ZN(_1455_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5025_ (.A1(_1430_),
    .A2(_1454_),
    .ZN(_1456_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5026_ (.A1(_1429_),
    .A2(_1456_),
    .ZN(_1457_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5027_ (.A1(_1418_),
    .A2(_1420_),
    .B(_1457_),
    .ZN(_1458_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5028_ (.A1(_1428_),
    .A2(_1457_),
    .ZN(_1459_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5029_ (.A1(_1427_),
    .A2(_1459_),
    .Z(_1460_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5030_ (.A1(_1241_),
    .A2(_1390_),
    .ZN(_1461_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5031_ (.A1(_1392_),
    .A2(_1461_),
    .Z(_1462_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5032_ (.A1(_1391_),
    .A2(_1460_),
    .B(_1462_),
    .ZN(_1463_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5033_ (.I(_1463_),
    .ZN(\dot2[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5034_ (.A1(_1427_),
    .A2(_1459_),
    .B(_1458_),
    .ZN(_1464_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5035_ (.A1(_1429_),
    .A2(_1456_),
    .B(_1455_),
    .ZN(_1465_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5036_ (.A1(net115),
    .A2(\pp_x_sq[10] ),
    .ZN(_1466_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5037_ (.A1(_1432_),
    .A2(_1453_),
    .B(_1452_),
    .ZN(_1467_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5038_ (.A1(_1401_),
    .A2(_1445_),
    .B1(_1447_),
    .B2(_1444_),
    .ZN(_1468_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5039_ (.I(_1468_),
    .ZN(_1469_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5040_ (.A1(_1441_),
    .A2(_1449_),
    .ZN(_1470_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5041_ (.A1(_1407_),
    .A2(_1436_),
    .B(_1439_),
    .ZN(_1471_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5042_ (.A1(net132),
    .A2(\pp_x_sq[14] ),
    .ZN(_1472_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5043_ (.A1(_1436_),
    .A2(_1472_),
    .Z(_1473_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5044_ (.A1(_1471_),
    .A2(_1473_),
    .ZN(_1474_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5045_ (.A1(_1471_),
    .A2(_1473_),
    .ZN(_1475_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5046_ (.I(_1475_),
    .ZN(_1476_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5047_ (.A1(net120),
    .A2(\pp_x_sq[11] ),
    .ZN(_1477_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5048_ (.A1(net124),
    .A2(\pp_x_sq[13] ),
    .ZN(_1478_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5049_ (.A1(net129),
    .A2(\pp_x_sq[13] ),
    .ZN(_1479_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5050_ (.A1(_1445_),
    .A2(_1479_),
    .ZN(_1480_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5051_ (.A1(_1477_),
    .A2(_1480_),
    .Z(_1481_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5052_ (.A1(_1476_),
    .A2(_1481_),
    .ZN(_1482_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5053_ (.A1(_1475_),
    .A2(_1481_),
    .Z(_1483_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5054_ (.I(_1483_),
    .ZN(_1484_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5055_ (.A1(_1470_),
    .A2(_1484_),
    .ZN(_1485_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5056_ (.A1(_1470_),
    .A2(_1484_),
    .ZN(_1486_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5057_ (.A1(_1468_),
    .A2(_1486_),
    .ZN(_1487_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5058_ (.A1(_1467_),
    .A2(_1487_),
    .ZN(_1488_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5059_ (.A1(_1467_),
    .A2(_1487_),
    .ZN(_1489_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5060_ (.A1(_1466_),
    .A2(_1489_),
    .ZN(_1490_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5061_ (.I(_1490_),
    .ZN(_1491_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5062_ (.A1(_1465_),
    .A2(_1491_),
    .ZN(_1492_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5063_ (.A1(_1465_),
    .A2(_1491_),
    .ZN(_1493_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5064_ (.A1(_1464_),
    .A2(_1465_),
    .A3(_1491_),
    .ZN(_1494_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5065_ (.A1(_1392_),
    .A2(_1494_),
    .ZN(_1495_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5066_ (.A1(_1240_),
    .A2(_1393_),
    .A3(_1425_),
    .ZN(_1496_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5067_ (.A1(_1391_),
    .A2(_1426_),
    .ZN(_1497_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5068_ (.A1(_1496_),
    .A2(_1497_),
    .B(_1495_),
    .ZN(\dot2[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5069_ (.A1(_1464_),
    .A2(_1493_),
    .B(_1492_),
    .ZN(_1498_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5070_ (.A1(_1466_),
    .A2(_1489_),
    .B(_1488_),
    .ZN(_1499_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5071_ (.I(_1499_),
    .ZN(_1500_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5072_ (.A1(net115),
    .A2(\pp_x_sq[11] ),
    .ZN(_1501_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5073_ (.A1(_1469_),
    .A2(_1486_),
    .B(_1485_),
    .ZN(_1502_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5074_ (.A1(_1446_),
    .A2(_1478_),
    .B1(_1480_),
    .B2(_1477_),
    .ZN(_1503_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5075_ (.I(_1503_),
    .ZN(_1504_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5076_ (.A1(_1474_),
    .A2(_1482_),
    .ZN(_1505_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5077_ (.A1(net132),
    .A2(\pp_x_sq[15] ),
    .A3(_1406_),
    .ZN(_1506_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5078_ (.A1(net120),
    .A2(\pp_x_sq[12] ),
    .ZN(_1507_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5079_ (.A1(net123),
    .A2(\pp_x_sq[14] ),
    .ZN(_1508_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5080_ (.A1(net129),
    .A2(\pp_x_sq[14] ),
    .ZN(_1509_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5081_ (.A1(_1478_),
    .A2(_1509_),
    .Z(_1510_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5082_ (.A1(net120),
    .A2(\pp_x_sq[12] ),
    .A3(_1510_),
    .ZN(_1511_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5083_ (.A1(_1507_),
    .A2(_1510_),
    .ZN(_1512_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _5084_ (.A1(net132),
    .A2(\pp_x_sq[15] ),
    .A3(_1406_),
    .A4(_1512_),
    .ZN(_1513_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5085_ (.A1(_1506_),
    .A2(_1512_),
    .ZN(_1514_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5086_ (.A1(_1505_),
    .A2(_1514_),
    .ZN(_1515_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5087_ (.A1(_1505_),
    .A2(_1514_),
    .ZN(_1516_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5088_ (.A1(_1503_),
    .A2(_1516_),
    .ZN(_1517_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5089_ (.A1(_1502_),
    .A2(_1517_),
    .ZN(_1518_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5090_ (.A1(_1502_),
    .A2(_1517_),
    .ZN(_1519_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5091_ (.A1(_1501_),
    .A2(_1519_),
    .ZN(_1520_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5092_ (.A1(_1500_),
    .A2(_1520_),
    .ZN(_1521_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5093_ (.A1(_1500_),
    .A2(_1520_),
    .ZN(_1522_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5094_ (.A1(_1498_),
    .A2(_1499_),
    .A3(_1520_),
    .ZN(_1523_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _5095_ (.I0(_1460_),
    .I1(_1523_),
    .S(_1392_),
    .Z(\dot2[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5096_ (.A1(_1498_),
    .A2(_1522_),
    .B(_1521_),
    .ZN(_1524_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5097_ (.A1(_1501_),
    .A2(_1519_),
    .B(_1518_),
    .ZN(_1525_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5098_ (.A1(net115),
    .A2(\pp_x_sq[12] ),
    .ZN(_1526_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5099_ (.A1(_1504_),
    .A2(_1516_),
    .B(_1515_),
    .ZN(_1527_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5100_ (.A1(_1479_),
    .A2(_1508_),
    .B(_1511_),
    .ZN(_1528_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5101_ (.I(_1528_),
    .ZN(_1529_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5102_ (.A1(_1436_),
    .A2(_1472_),
    .B(_1513_),
    .ZN(_1530_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5103_ (.A1(net129),
    .A2(\pp_x_sq[15] ),
    .ZN(_1531_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5104_ (.A1(net123),
    .A2(\pp_x_sq[15] ),
    .ZN(_1532_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5105_ (.A1(_1508_),
    .A2(_1531_),
    .Z(_1533_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5106_ (.A1(net120),
    .A2(\pp_x_sq[13] ),
    .ZN(_1534_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5107_ (.A1(net120),
    .A2(\pp_x_sq[13] ),
    .A3(_1533_),
    .ZN(_1535_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5108_ (.A1(_1533_),
    .A2(_1534_),
    .ZN(_1536_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5109_ (.A1(_1530_),
    .A2(_1536_),
    .ZN(_1537_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5110_ (.A1(_1529_),
    .A2(_1537_),
    .ZN(_1538_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5111_ (.A1(_1528_),
    .A2(_1537_),
    .ZN(_1539_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5112_ (.A1(_1527_),
    .A2(_1539_),
    .ZN(_1540_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5113_ (.A1(_1527_),
    .A2(_1539_),
    .ZN(_1541_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5114_ (.A1(_1526_),
    .A2(_1541_),
    .ZN(_1542_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5115_ (.I(_1542_),
    .ZN(_1543_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5116_ (.A1(_1525_),
    .A2(_1543_),
    .ZN(_1544_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5117_ (.A1(_1525_),
    .A2(_1543_),
    .ZN(_1545_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5118_ (.A1(_1524_),
    .A2(_1525_),
    .A3(_1543_),
    .ZN(_1546_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _5119_ (.I0(_1494_),
    .I1(_1546_),
    .S(_1392_),
    .Z(\dot2[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5120_ (.A1(_1524_),
    .A2(_1545_),
    .B(_1544_),
    .ZN(_1547_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5121_ (.A1(_1526_),
    .A2(_1541_),
    .B(_1540_),
    .ZN(_1548_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5122_ (.I(_1548_),
    .ZN(_1549_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5123_ (.A1(net115),
    .A2(\pp_x_sq[13] ),
    .ZN(_1550_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5124_ (.A1(net121),
    .A2(\pp_x_sq[14] ),
    .ZN(_1551_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5125_ (.A1(_1532_),
    .A2(_1551_),
    .Z(_1552_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5126_ (.A1(_1532_),
    .A2(_1551_),
    .Z(_1553_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5127_ (.A1(_1509_),
    .A2(_1532_),
    .B(_1535_),
    .ZN(_1554_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5128_ (.A1(_1553_),
    .A2(_1554_),
    .ZN(_1555_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5129_ (.A1(_1553_),
    .A2(_1554_),
    .ZN(_1556_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5130_ (.A1(_1530_),
    .A2(_1536_),
    .B(_1538_),
    .ZN(_1557_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5131_ (.A1(_1556_),
    .A2(_1557_),
    .Z(_1558_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5132_ (.A1(_1556_),
    .A2(_1557_),
    .ZN(_1559_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5133_ (.A1(_1558_),
    .A2(_1559_),
    .ZN(_1560_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5134_ (.A1(_1550_),
    .A2(_1560_),
    .ZN(_1561_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5135_ (.A1(_1549_),
    .A2(_1561_),
    .ZN(_1562_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5136_ (.A1(_1549_),
    .A2(_1561_),
    .ZN(_1563_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5137_ (.A1(_1547_),
    .A2(_1548_),
    .A3(_1561_),
    .ZN(_1564_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _5138_ (.I0(_1523_),
    .I1(_1564_),
    .S(_1392_),
    .Z(\dot2[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5139_ (.A1(_1547_),
    .A2(_1563_),
    .B(_1562_),
    .ZN(_1565_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5140_ (.A1(_1550_),
    .A2(_1560_),
    .B(_1558_),
    .ZN(_1566_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5141_ (.A1(net113),
    .A2(\pp_x_sq[14] ),
    .ZN(_1567_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5142_ (.A1(net121),
    .A2(\pp_x_sq[15] ),
    .A3(_1508_),
    .ZN(_1568_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5143_ (.A1(_1555_),
    .A2(_1568_),
    .ZN(_1569_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5144_ (.A1(_1555_),
    .A2(_1568_),
    .ZN(_1570_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5145_ (.A1(_1567_),
    .A2(_1570_),
    .ZN(_1571_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5146_ (.A1(_1567_),
    .A2(_1570_),
    .Z(_1572_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5147_ (.A1(_1566_),
    .A2(_1572_),
    .ZN(_1573_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5148_ (.A1(_1566_),
    .A2(_1572_),
    .ZN(_1574_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5149_ (.A1(_1565_),
    .A2(_1566_),
    .A3(_1572_),
    .ZN(_1575_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _5150_ (.I0(_1546_),
    .I1(_1575_),
    .S(_1392_),
    .Z(\dot2[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5151_ (.A1(net113),
    .A2(\pp_x_sq[15] ),
    .ZN(_1576_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _5152_ (.I0(net113),
    .I1(_1576_),
    .S(_1552_),
    .Z(_1577_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5153_ (.A1(_1569_),
    .A2(_1571_),
    .ZN(_1578_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5154_ (.A1(_1577_),
    .A2(_1578_),
    .Z(_1579_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5155_ (.A1(_1577_),
    .A2(_1578_),
    .ZN(_1580_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5156_ (.A1(_1579_),
    .A2(_1580_),
    .ZN(_1581_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5157_ (.A1(_1565_),
    .A2(_1574_),
    .B(_1573_),
    .ZN(_1582_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5158_ (.A1(_1581_),
    .A2(_1582_),
    .ZN(_1583_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _5159_ (.I0(_1564_),
    .I1(_1583_),
    .S(_1392_),
    .Z(\dot2[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5160_ (.A1(_1580_),
    .A2(_1582_),
    .ZN(_1584_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5161_ (.A1(net88),
    .A2(_1552_),
    .B(_1579_),
    .C(_1584_),
    .ZN(_1585_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _5162_ (.I0(_1575_),
    .I1(_1585_),
    .S(_1392_),
    .Z(\dot2[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _5163_ (.A1(net113),
    .A2(_0081_),
    .A3(_2773_),
    .A4(_2776_),
    .ZN(_0012_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5164_ (.A1(_2704_),
    .A2(_2706_),
    .B(_2701_),
    .ZN(_1586_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _5165_ (.A1(net116),
    .A2(_2571_),
    .B(_2720_),
    .C(_1586_),
    .ZN(_1587_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_1 _5166_ (.A1(net153),
    .A2(_2627_),
    .A3(_2719_),
    .A4(_1587_),
    .ZN(_1588_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _5167_ (.A1(net154),
    .A2(_2627_),
    .A3(_2719_),
    .A4(_1587_),
    .Z(_1589_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5168_ (.A1(net136),
    .A2(\r2[0] ),
    .ZN(_1590_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5169_ (.A1(net136),
    .A2(\r2[0] ),
    .ZN(_1591_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _5170_ (.A1(_2573_),
    .A2(_2576_),
    .B(_2575_),
    .ZN(_1592_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5171_ (.A1(\hvsync_gen.hpos[9] ),
    .A2(_2746_),
    .ZN(_1593_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5172_ (.A1(net62),
    .A2(_2752_),
    .ZN(_1594_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5173_ (.A1(net76),
    .A2(_2751_),
    .ZN(_1595_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _5174_ (.A1(_1593_),
    .A2(net47),
    .ZN(_1596_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5175_ (.A1(_1592_),
    .A2(net46),
    .ZN(_1597_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5176_ (.A1(\r2[0] ),
    .A2(net84),
    .Z(_1598_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5177_ (.A1(net22),
    .A2(_1598_),
    .ZN(_1599_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5178_ (.A1(net22),
    .A2(_1591_),
    .B(net42),
    .C(_1599_),
    .ZN(_1600_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5179_ (.A1(_2760_),
    .A2(_1592_),
    .ZN(_1601_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5180_ (.A1(_2760_),
    .A2(_1592_),
    .Z(_1602_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _5181_ (.A1(net47),
    .A2(net37),
    .ZN(_1603_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5182_ (.A1(net46),
    .A2(net33),
    .ZN(_1604_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and4_1 _5183_ (.A1(\hvsync_gen.vpos[5] ),
    .A2(net92),
    .A3(\hvsync_gen.vpos[7] ),
    .A4(\hvsync_gen.vpos[8] ),
    .Z(_1605_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _5184_ (.A1(\hvsync_gen.vpos[9] ),
    .A2(_1605_),
    .ZN(_1606_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5185_ (.A1(_1593_),
    .A2(_1606_),
    .Z(_1607_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5186_ (.A1(_1593_),
    .A2(_1606_),
    .ZN(_1608_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5187_ (.A1(net59),
    .A2(_1608_),
    .ZN(_1609_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5188_ (.A1(net58),
    .A2(_1607_),
    .ZN(_1610_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5189_ (.A1(_1598_),
    .A2(net30),
    .ZN(_1611_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5190_ (.A1(\r2[0] ),
    .A2(net30),
    .B(_1611_),
    .C(net40),
    .ZN(_1612_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5191_ (.A1(_1600_),
    .A2(net21),
    .A3(_1612_),
    .ZN(_1613_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5192_ (.A1(_1598_),
    .A2(net39),
    .ZN(_1614_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5193_ (.A1(_1613_),
    .A2(_1614_),
    .B(net165),
    .ZN(_0013_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5194_ (.A1(net131),
    .A2(\r2[1] ),
    .ZN(_1615_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5195_ (.A1(net131),
    .A2(\r2[1] ),
    .ZN(_1616_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5196_ (.A1(_2550_),
    .A2(_2597_),
    .A3(_1590_),
    .ZN(_1617_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5197_ (.A1(net23),
    .A2(_1617_),
    .ZN(_1618_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5198_ (.A1(net89),
    .A2(_2597_),
    .ZN(_1619_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5199_ (.A1(_1589_),
    .A2(_1619_),
    .B(net41),
    .ZN(_1620_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5200_ (.A1(\r2[1] ),
    .A2(_2630_),
    .ZN(_1621_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5201_ (.A1(\r2[0] ),
    .A2(_1621_),
    .Z(_1622_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5202_ (.A1(\r2[0] ),
    .A2(_1621_),
    .ZN(_1623_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5203_ (.A1(net32),
    .A2(_1622_),
    .A3(_1623_),
    .ZN(_1624_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5204_ (.A1(net30),
    .A2(_1619_),
    .B(net42),
    .ZN(_1625_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5205_ (.A1(_1618_),
    .A2(_1620_),
    .B1(_1624_),
    .B2(_1625_),
    .ZN(_1626_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5206_ (.A1(net39),
    .A2(_1619_),
    .B1(_1626_),
    .B2(_1603_),
    .ZN(_1627_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5207_ (.A1(net166),
    .A2(_1627_),
    .ZN(_0014_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5208_ (.A1(net89),
    .A2(_2598_),
    .ZN(_1628_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5209_ (.A1(_1590_),
    .A2(_1616_),
    .B(_1615_),
    .ZN(_1629_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5210_ (.A1(net126),
    .A2(\r2[2] ),
    .ZN(_1630_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5211_ (.A1(net126),
    .A2(\r2[2] ),
    .Z(_1631_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5212_ (.A1(_1629_),
    .A2(_1631_),
    .ZN(_1632_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5213_ (.A1(_1629_),
    .A2(_1631_),
    .ZN(_1633_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5214_ (.A1(_2597_),
    .A2(_2630_),
    .B(_1623_),
    .ZN(_1634_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5215_ (.A1(_2598_),
    .A2(_2653_),
    .ZN(_1635_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5216_ (.A1(_2598_),
    .A2(_2653_),
    .ZN(_1636_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5217_ (.A1(net24),
    .A2(_1633_),
    .ZN(_1637_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5218_ (.A1(net24),
    .A2(_1628_),
    .B(_1637_),
    .C(net42),
    .ZN(_1638_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5219_ (.A1(_2598_),
    .A2(_2653_),
    .A3(_1634_),
    .ZN(_1639_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5220_ (.A1(net32),
    .A2(_1639_),
    .ZN(_1640_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5221_ (.A1(net32),
    .A2(_1628_),
    .B(_1640_),
    .C(net41),
    .ZN(_1641_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5222_ (.A1(_1638_),
    .A2(_1641_),
    .ZN(_1642_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5223_ (.A1(net39),
    .A2(_1628_),
    .B1(_1642_),
    .B2(net21),
    .ZN(_1643_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5224_ (.A1(net166),
    .A2(_1643_),
    .ZN(_0015_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5225_ (.A1(net90),
    .A2(_2599_),
    .ZN(_1644_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5226_ (.A1(_1630_),
    .A2(_1632_),
    .ZN(_1645_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5227_ (.A1(_2548_),
    .A2(_2599_),
    .ZN(_1646_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5228_ (.A1(net123),
    .A2(\r2[3] ),
    .ZN(_1647_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5229_ (.A1(_1630_),
    .A2(_1632_),
    .B(_1647_),
    .ZN(_1648_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5230_ (.A1(_1645_),
    .A2(_1647_),
    .Z(_1649_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5231_ (.A1(net24),
    .A2(_1649_),
    .ZN(_1650_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5232_ (.A1(net24),
    .A2(_1644_),
    .B(_1650_),
    .C(net42),
    .ZN(_1651_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5233_ (.A1(_1634_),
    .A2(_1636_),
    .B(_1635_),
    .ZN(_1652_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5234_ (.A1(\r2[3] ),
    .A2(_2667_),
    .A3(_2668_),
    .ZN(_1653_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5235_ (.A1(_2599_),
    .A2(_2669_),
    .ZN(_1654_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5236_ (.A1(net32),
    .A2(_1644_),
    .ZN(_1655_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5237_ (.A1(_1652_),
    .A2(_1654_),
    .Z(_1656_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5238_ (.A1(net30),
    .A2(_1656_),
    .ZN(_1657_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _5239_ (.A1(net42),
    .A2(_1655_),
    .A3(_1657_),
    .B(_1651_),
    .ZN(_1658_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5240_ (.A1(net38),
    .A2(_1644_),
    .B1(_1658_),
    .B2(_1603_),
    .ZN(_1659_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5241_ (.A1(net168),
    .A2(_1659_),
    .ZN(_0016_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5242_ (.A1(_2600_),
    .A2(_2686_),
    .ZN(_1660_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5243_ (.A1(\r2[4] ),
    .A2(_2686_),
    .ZN(_1661_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _5244_ (.A1(_1652_),
    .A2(_1654_),
    .B(_1653_),
    .ZN(_1662_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5245_ (.A1(_1661_),
    .A2(_1662_),
    .ZN(_1663_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5246_ (.A1(_1661_),
    .A2(_1662_),
    .ZN(_1664_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5247_ (.A1(net30),
    .A2(_1663_),
    .ZN(_1665_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5248_ (.A1(net90),
    .A2(_2600_),
    .ZN(_1666_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5249_ (.A1(_1664_),
    .A2(_1665_),
    .B1(_1666_),
    .B2(net31),
    .C(_1596_),
    .ZN(_1667_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5250_ (.A1(net86),
    .A2(_2600_),
    .ZN(_1668_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5251_ (.A1(net86),
    .A2(_2600_),
    .ZN(_1669_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5252_ (.A1(_1646_),
    .A2(_1648_),
    .Z(_1670_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5253_ (.A1(net121),
    .A2(_2600_),
    .A3(_1670_),
    .ZN(_1671_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5254_ (.A1(net24),
    .A2(_1671_),
    .ZN(_1672_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5255_ (.A1(_1589_),
    .A2(_1666_),
    .B(net41),
    .ZN(_1673_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _5256_ (.A1(_1672_),
    .A2(_1673_),
    .B(_1604_),
    .C(_1667_),
    .ZN(_1674_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5257_ (.A1(net38),
    .A2(_1666_),
    .B(_1674_),
    .ZN(_1675_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5258_ (.A1(net166),
    .A2(_1675_),
    .ZN(_0017_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5259_ (.A1(net90),
    .A2(_2601_),
    .ZN(_1676_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5260_ (.A1(net112),
    .A2(\r2[5] ),
    .ZN(_1677_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5261_ (.A1(net112),
    .A2(\r2[5] ),
    .ZN(_1678_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5262_ (.A1(_1669_),
    .A2(_1670_),
    .B(_1668_),
    .ZN(_1679_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5263_ (.A1(net88),
    .A2(\r2[5] ),
    .A3(_1679_),
    .ZN(_1680_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5264_ (.A1(net24),
    .A2(_1680_),
    .ZN(_1681_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5265_ (.A1(net24),
    .A2(_1676_),
    .B(_1681_),
    .C(_1596_),
    .ZN(_1682_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5266_ (.A1(_1661_),
    .A2(_1662_),
    .B(_1660_),
    .ZN(_1683_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5267_ (.A1(\r2[5] ),
    .A2(_2708_),
    .ZN(_1684_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5268_ (.A1(_2601_),
    .A2(_2708_),
    .A3(_1683_),
    .ZN(_1685_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5269_ (.A1(net32),
    .A2(_1685_),
    .ZN(_1686_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5270_ (.A1(net32),
    .A2(_1676_),
    .B(_1686_),
    .C(net41),
    .ZN(_1687_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5271_ (.A1(_1682_),
    .A2(_1687_),
    .ZN(_1688_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5272_ (.A1(net38),
    .A2(_1676_),
    .B1(_1688_),
    .B2(_1603_),
    .ZN(_1689_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5273_ (.A1(net166),
    .A2(_1689_),
    .ZN(_0018_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5274_ (.A1(\r2[6] ),
    .A2(_2723_),
    .ZN(_1690_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5275_ (.A1(\r2[6] ),
    .A2(_2723_),
    .ZN(_1691_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _5276_ (.A1(\r2[5] ),
    .A2(_2708_),
    .B1(_1661_),
    .B2(_1662_),
    .C(_1660_),
    .ZN(_1692_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5277_ (.A1(_1684_),
    .A2(_1692_),
    .Z(_1693_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5278_ (.A1(_1691_),
    .A2(_1693_),
    .ZN(_1694_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5279_ (.A1(net58),
    .A2(_1606_),
    .A3(_1694_),
    .ZN(_1695_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5280_ (.A1(net83),
    .A2(\r2[6] ),
    .ZN(_1696_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5281_ (.A1(_1592_),
    .A2(_1696_),
    .B(net30),
    .ZN(_1697_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5282_ (.A1(_2760_),
    .A2(_1695_),
    .A3(_1697_),
    .ZN(_1698_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5283_ (.A1(_1678_),
    .A2(_1679_),
    .B(_1677_),
    .ZN(_1699_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5284_ (.A1(net24),
    .A2(_1699_),
    .ZN(_1700_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5285_ (.A1(\r2[6] ),
    .A2(_1699_),
    .ZN(_1701_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5286_ (.A1(net89),
    .A2(net22),
    .ZN(_1702_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5287_ (.A1(net42),
    .A2(_1702_),
    .ZN(_1703_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5288_ (.A1(\r2[6] ),
    .A2(_1700_),
    .Z(_1704_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai221_1 _5289_ (.A1(net33),
    .A2(_1696_),
    .B1(_1703_),
    .B2(_1704_),
    .C(_1698_),
    .ZN(_1705_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5290_ (.A1(net169),
    .A2(_1705_),
    .Z(_0019_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5291_ (.A1(net84),
    .A2(\r2[7] ),
    .ZN(_1706_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5292_ (.A1(\r2[7] ),
    .A2(_2735_),
    .ZN(_1707_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5293_ (.A1(_2602_),
    .A2(_2735_),
    .ZN(_1708_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _5294_ (.A1(_1684_),
    .A2(_1691_),
    .A3(_1692_),
    .B(_1690_),
    .ZN(_1709_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5295_ (.A1(_1708_),
    .A2(_1709_),
    .ZN(_1710_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5296_ (.A1(_1708_),
    .A2(_1709_),
    .Z(_1711_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5297_ (.A1(net41),
    .A2(net30),
    .A3(_1706_),
    .ZN(_1712_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5298_ (.A1(_1603_),
    .A2(_1712_),
    .ZN(_1713_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5299_ (.A1(_2602_),
    .A2(_1701_),
    .B(_1589_),
    .ZN(_1714_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5300_ (.A1(\r2[6] ),
    .A2(\r2[7] ),
    .A3(_1699_),
    .ZN(_1715_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5301_ (.A1(_1589_),
    .A2(_1706_),
    .B1(_1714_),
    .B2(_1715_),
    .ZN(_1716_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5302_ (.A1(net30),
    .A2(_1711_),
    .B1(_1716_),
    .B2(net41),
    .ZN(_1717_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5303_ (.A1(net34),
    .A2(_1706_),
    .B1(_1713_),
    .B2(_1717_),
    .ZN(_1718_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5304_ (.A1(net169),
    .A2(_1718_),
    .Z(_0020_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5305_ (.A1(net84),
    .A2(\r2[8] ),
    .A3(net38),
    .ZN(_1719_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5306_ (.A1(_1707_),
    .A2(_1710_),
    .ZN(_1720_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5307_ (.A1(_0462_),
    .A2(_0463_),
    .B(_2603_),
    .ZN(_1721_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5308_ (.A1(\r2[8] ),
    .A2(_0464_),
    .ZN(_1722_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5309_ (.A1(_1707_),
    .A2(_1710_),
    .B(_1722_),
    .ZN(_1723_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5310_ (.A1(_1720_),
    .A2(_1722_),
    .Z(_1724_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5311_ (.A1(net84),
    .A2(\r2[8] ),
    .B(_1609_),
    .ZN(_1725_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _5312_ (.A1(_1609_),
    .A2(_1724_),
    .B(_1725_),
    .C(_1596_),
    .ZN(_1726_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5313_ (.A1(\r2[8] ),
    .A2(_1714_),
    .ZN(_1727_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5314_ (.A1(_1703_),
    .A2(_1727_),
    .ZN(_1728_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5315_ (.A1(_1726_),
    .A2(_1728_),
    .B(net21),
    .ZN(_1729_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5316_ (.A1(_1719_),
    .A2(_1729_),
    .B(net165),
    .ZN(_0021_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5317_ (.A1(net82),
    .A2(\r2[9] ),
    .A3(net37),
    .ZN(_1730_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5318_ (.A1(\r2[9] ),
    .A2(_0533_),
    .Z(_1731_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5319_ (.A1(\r2[9] ),
    .A2(_0533_),
    .Z(_1732_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5320_ (.A1(_1721_),
    .A2(_1732_),
    .Z(_1733_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _5321_ (.A1(_1723_),
    .A2(_1732_),
    .B(_1733_),
    .C(net30),
    .ZN(_1734_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _5322_ (.A1(_1721_),
    .A2(_1723_),
    .A3(_1732_),
    .B(_1734_),
    .ZN(_1735_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5323_ (.A1(net83),
    .A2(\r2[9] ),
    .A3(net30),
    .ZN(_1736_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5324_ (.A1(net40),
    .A2(_1735_),
    .A3(_1736_),
    .ZN(_1737_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5325_ (.A1(_2602_),
    .A2(_1701_),
    .B(_2603_),
    .ZN(_1738_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5326_ (.A1(\r2[9] ),
    .A2(net22),
    .A3(_1738_),
    .ZN(_1739_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5327_ (.A1(net22),
    .A2(_1738_),
    .B(_1702_),
    .C(\r2[9] ),
    .ZN(_1740_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5328_ (.A1(_1592_),
    .A2(_1740_),
    .ZN(_1741_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5329_ (.A1(_1739_),
    .A2(_1741_),
    .B(net21),
    .C(_1737_),
    .ZN(_1742_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5330_ (.A1(_1730_),
    .A2(_1742_),
    .B(net165),
    .ZN(_0022_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5331_ (.A1(net89),
    .A2(_2604_),
    .ZN(_1743_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5332_ (.A1(_2575_),
    .A2(_0532_),
    .ZN(_1744_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5333_ (.A1(\r2[10] ),
    .A2(net15),
    .ZN(_1745_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5334_ (.A1(\r2[10] ),
    .A2(net15),
    .ZN(_1746_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _5335_ (.A1(_1723_),
    .A2(_1732_),
    .B(_1733_),
    .C(_1731_),
    .ZN(_1747_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5336_ (.A1(_2604_),
    .A2(net15),
    .A3(_1747_),
    .ZN(_1748_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5337_ (.A1(net32),
    .A2(_1748_),
    .ZN(_1749_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5338_ (.A1(net32),
    .A2(_1743_),
    .B(_1749_),
    .C(net40),
    .ZN(_1750_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5339_ (.A1(\r2[9] ),
    .A2(_1738_),
    .ZN(_1751_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5340_ (.A1(net22),
    .A2(_1751_),
    .ZN(_1752_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5341_ (.A1(\r2[10] ),
    .A2(_1752_),
    .ZN(_1753_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5342_ (.A1(_1703_),
    .A2(_1753_),
    .B(_1750_),
    .ZN(_1754_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5343_ (.A1(net37),
    .A2(_1743_),
    .B1(_1754_),
    .B2(net21),
    .ZN(_1755_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5344_ (.A1(net165),
    .A2(_1755_),
    .ZN(_0023_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5345_ (.A1(_1746_),
    .A2(_1747_),
    .B(_1745_),
    .ZN(_1756_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5346_ (.A1(\r2[11] ),
    .A2(net15),
    .ZN(_1757_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _5347_ (.A1(\r2[11] ),
    .A2(net15),
    .A3(_1756_),
    .Z(_1758_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5348_ (.A1(_2754_),
    .A2(_1608_),
    .ZN(_1759_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5349_ (.A1(net59),
    .A2(_1606_),
    .ZN(_1760_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5350_ (.A1(net82),
    .A2(\r2[11] ),
    .ZN(_1761_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5351_ (.A1(_1608_),
    .A2(_1761_),
    .ZN(_1762_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5352_ (.A1(_1608_),
    .A2(_1758_),
    .B(net44),
    .C(_1762_),
    .ZN(_1763_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5353_ (.A1(net44),
    .A2(_1761_),
    .B(_1763_),
    .C(net40),
    .ZN(_1764_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5354_ (.A1(_2604_),
    .A2(_1751_),
    .ZN(_1765_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5355_ (.A1(\r2[11] ),
    .A2(_1765_),
    .ZN(_1766_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5356_ (.A1(\r2[11] ),
    .A2(_1765_),
    .ZN(_1767_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5357_ (.A1(net23),
    .A2(_1766_),
    .ZN(_1768_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5358_ (.A1(net23),
    .A2(_1761_),
    .B1(_1767_),
    .B2(_1768_),
    .ZN(_1769_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5359_ (.A1(net40),
    .A2(_1769_),
    .B(_1764_),
    .ZN(_1770_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5360_ (.A1(net33),
    .A2(_1761_),
    .B1(_1770_),
    .B2(_1604_),
    .ZN(_1771_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5361_ (.A1(net170),
    .A2(_1771_),
    .Z(_0024_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5362_ (.A1(_2605_),
    .A2(net14),
    .ZN(_1772_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5363_ (.I(_1772_),
    .ZN(_1773_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5364_ (.A1(\r2[11] ),
    .A2(net14),
    .B(_1756_),
    .ZN(_1774_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5365_ (.A1(_1757_),
    .A2(_1774_),
    .ZN(_1775_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5366_ (.A1(_1757_),
    .A2(_1774_),
    .B(_1773_),
    .ZN(_1776_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5367_ (.A1(net31),
    .A2(_1776_),
    .ZN(_1777_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5368_ (.A1(_1772_),
    .A2(_1775_),
    .B(_1777_),
    .ZN(_1778_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5369_ (.A1(_2605_),
    .A2(_1766_),
    .ZN(_1779_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5370_ (.A1(\r2[11] ),
    .A2(_1765_),
    .B(\r2[12] ),
    .ZN(_1780_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5371_ (.A1(_1779_),
    .A2(_1780_),
    .B(net23),
    .ZN(_1781_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5372_ (.A1(net83),
    .A2(\r2[12] ),
    .ZN(_1782_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5373_ (.A1(net22),
    .A2(_1782_),
    .B(_1593_),
    .ZN(_1783_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _5374_ (.A1(_1592_),
    .A2(net32),
    .A3(_1782_),
    .B(net21),
    .ZN(_1784_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5375_ (.A1(_1781_),
    .A2(_1783_),
    .B(_1784_),
    .ZN(_1785_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5376_ (.A1(net37),
    .A2(_1782_),
    .B1(_1785_),
    .B2(_1778_),
    .C(net167),
    .ZN(_0025_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5377_ (.A1(net83),
    .A2(\r2[13] ),
    .ZN(_1786_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5378_ (.A1(net83),
    .A2(\r2[13] ),
    .A3(net37),
    .ZN(_1787_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5379_ (.A1(_2606_),
    .A2(net14),
    .ZN(_1788_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5380_ (.A1(\r2[12] ),
    .A2(net14),
    .B(_1776_),
    .ZN(_1789_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5381_ (.A1(_1788_),
    .A2(_1789_),
    .B(_1608_),
    .ZN(_1790_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5382_ (.A1(_1788_),
    .A2(_1789_),
    .B(_1790_),
    .ZN(_1791_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5383_ (.A1(_1608_),
    .A2(_1786_),
    .ZN(_1792_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5384_ (.A1(net44),
    .A2(_1791_),
    .A3(_1792_),
    .ZN(_1793_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5385_ (.A1(net44),
    .A2(_1786_),
    .B(_1793_),
    .C(net40),
    .ZN(_1794_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5386_ (.A1(_2605_),
    .A2(_2606_),
    .A3(_1766_),
    .ZN(_1795_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5387_ (.A1(\r2[13] ),
    .A2(_1779_),
    .B(net23),
    .ZN(_1796_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5388_ (.A1(net23),
    .A2(_1786_),
    .B1(_1795_),
    .B2(_1796_),
    .ZN(_1797_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5389_ (.A1(net40),
    .A2(_1797_),
    .B(_1794_),
    .C(net21),
    .ZN(_1798_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5390_ (.A1(_1787_),
    .A2(_1798_),
    .B(net165),
    .ZN(_0026_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5391_ (.A1(\r2[14] ),
    .A2(net14),
    .ZN(_1799_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5392_ (.A1(_2607_),
    .A2(net14),
    .ZN(_1800_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5393_ (.A1(_1776_),
    .A2(_1788_),
    .ZN(_1801_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5394_ (.A1(\r2[12] ),
    .A2(\r2[13] ),
    .B(net15),
    .ZN(_1802_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5395_ (.A1(_1801_),
    .A2(_1802_),
    .ZN(_1803_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5396_ (.A1(_1800_),
    .A2(_1803_),
    .ZN(_1804_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5397_ (.A1(_1800_),
    .A2(_1803_),
    .ZN(_1805_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5398_ (.A1(net32),
    .A2(_1805_),
    .ZN(_1806_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5399_ (.A1(\r2[14] ),
    .A2(_1795_),
    .Z(_1807_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5400_ (.A1(\r2[14] ),
    .A2(_1795_),
    .B(net23),
    .ZN(_1808_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5401_ (.A1(net82),
    .A2(\r2[14] ),
    .ZN(_1809_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai221_1 _5402_ (.A1(_1807_),
    .A2(_1808_),
    .B1(_1809_),
    .B2(net23),
    .C(net42),
    .ZN(_1810_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5403_ (.A1(net40),
    .A2(net31),
    .A3(_1809_),
    .ZN(_1811_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _5404_ (.A1(net21),
    .A2(_1806_),
    .A3(_1810_),
    .A4(_1811_),
    .ZN(_1812_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5405_ (.A1(net82),
    .A2(\r2[14] ),
    .A3(net35),
    .ZN(_1813_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5406_ (.A1(_1812_),
    .A2(_1813_),
    .B(net164),
    .ZN(_0027_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5407_ (.A1(\r2[15] ),
    .A2(net14),
    .ZN(_1814_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5408_ (.A1(\r2[15] ),
    .A2(net14),
    .Z(_1815_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5409_ (.A1(_1799_),
    .A2(_1804_),
    .A3(_1815_),
    .ZN(_1816_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5410_ (.A1(_1799_),
    .A2(_1804_),
    .B(_1815_),
    .ZN(_1817_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5411_ (.A1(net31),
    .A2(_1817_),
    .ZN(_1818_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5412_ (.A1(_1816_),
    .A2(_1818_),
    .ZN(_1819_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5413_ (.A1(net82),
    .A2(\r2[15] ),
    .ZN(_1820_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5414_ (.A1(net31),
    .A2(_1820_),
    .B(net42),
    .ZN(_1821_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5415_ (.A1(net23),
    .A2(_1807_),
    .B(\r2[15] ),
    .ZN(_1822_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5416_ (.A1(\r2[15] ),
    .A2(net23),
    .A3(_1807_),
    .ZN(_1823_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5417_ (.A1(_1592_),
    .A2(_1702_),
    .A3(_1823_),
    .ZN(_1824_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5418_ (.A1(_1822_),
    .A2(_1824_),
    .B(net21),
    .ZN(_1825_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5419_ (.A1(_1819_),
    .A2(_1821_),
    .B(_1825_),
    .ZN(_1826_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _5420_ (.A1(net37),
    .A2(_1820_),
    .B(_1826_),
    .C(net165),
    .ZN(_0028_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5421_ (.A1(\r2[16] ),
    .A2(net15),
    .ZN(_1827_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5422_ (.A1(\r2[16] ),
    .A2(net14),
    .Z(_1828_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and4_1 _5423_ (.A1(_1776_),
    .A2(_1788_),
    .A3(_1800_),
    .A4(_1815_),
    .Z(_1829_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5424_ (.A1(_1799_),
    .A2(_1802_),
    .A3(_1814_),
    .ZN(_1830_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5425_ (.A1(_1829_),
    .A2(_1830_),
    .ZN(_1831_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5426_ (.A1(_1829_),
    .A2(_1830_),
    .B(_1828_),
    .ZN(_1832_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5427_ (.A1(_1828_),
    .A2(_1831_),
    .ZN(_1833_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5428_ (.A1(\r2[16] ),
    .A2(_1702_),
    .A3(_1823_),
    .ZN(_1834_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5429_ (.A1(\r2[16] ),
    .A2(_1823_),
    .B(_1834_),
    .C(net42),
    .ZN(_1835_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5430_ (.A1(net82),
    .A2(\r2[16] ),
    .ZN(_1836_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5431_ (.A1(_1593_),
    .A2(net31),
    .A3(_1836_),
    .ZN(_1837_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5432_ (.A1(net31),
    .A2(_1833_),
    .B(_1835_),
    .C(_1837_),
    .ZN(_1838_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5433_ (.A1(net37),
    .A2(_1836_),
    .ZN(_1839_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5434_ (.A1(net170),
    .A2(_1839_),
    .ZN(_1840_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5435_ (.A1(net33),
    .A2(_1838_),
    .B(_1840_),
    .ZN(_0029_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5436_ (.A1(net89),
    .A2(_2608_),
    .ZN(_1841_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5437_ (.A1(net37),
    .A2(_1841_),
    .ZN(_1842_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5438_ (.A1(_1827_),
    .A2(_1832_),
    .ZN(_1843_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5439_ (.A1(\r2[17] ),
    .A2(net15),
    .ZN(_1844_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5440_ (.A1(_1827_),
    .A2(_1832_),
    .A3(_1844_),
    .ZN(_1845_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5441_ (.A1(_2608_),
    .A2(_1744_),
    .A3(_1843_),
    .ZN(_1846_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5442_ (.A1(_1608_),
    .A2(_1846_),
    .ZN(_1847_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5443_ (.A1(_1607_),
    .A2(_1841_),
    .B(net45),
    .ZN(_1848_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5444_ (.A1(net28),
    .A2(_1841_),
    .ZN(_1849_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5445_ (.A1(_1847_),
    .A2(_1848_),
    .B(_1849_),
    .C(net40),
    .ZN(_1850_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5446_ (.A1(\r2[15] ),
    .A2(\r2[16] ),
    .A3(_1807_),
    .ZN(_1851_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5447_ (.A1(_2608_),
    .A2(_1851_),
    .ZN(_1852_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5448_ (.A1(net22),
    .A2(_1841_),
    .ZN(_1853_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5449_ (.A1(net22),
    .A2(_1852_),
    .B(_1853_),
    .C(net42),
    .ZN(_1854_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5450_ (.A1(net21),
    .A2(_1850_),
    .A3(_1854_),
    .ZN(_1855_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5451_ (.A1(_1842_),
    .A2(_1855_),
    .B(net165),
    .ZN(_0030_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5452_ (.A1(\r2[17] ),
    .A2(net15),
    .B(_1845_),
    .ZN(_1856_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5453_ (.A1(\r2[18] ),
    .A2(net14),
    .A3(_1856_),
    .ZN(_1857_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or3_1 _5454_ (.A1(_2608_),
    .A2(net22),
    .A3(_1851_),
    .Z(_1858_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5455_ (.A1(\r2[18] ),
    .A2(_1702_),
    .ZN(_1859_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _5456_ (.I0(\r2[18] ),
    .I1(_1859_),
    .S(_1858_),
    .Z(_1860_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5457_ (.A1(net82),
    .A2(\r2[18] ),
    .ZN(_1861_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5458_ (.A1(net40),
    .A2(net31),
    .A3(_1861_),
    .ZN(_1862_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5459_ (.A1(_1592_),
    .A2(_1860_),
    .B(_1604_),
    .ZN(_1863_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5460_ (.A1(net31),
    .A2(_1857_),
    .B(_1862_),
    .C(_1863_),
    .ZN(_1864_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5461_ (.A1(net82),
    .A2(\r2[18] ),
    .A3(net35),
    .ZN(_1865_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5462_ (.A1(_1864_),
    .A2(_1865_),
    .B(net164),
    .ZN(_0031_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5463_ (.A1(net113),
    .A2(_0081_),
    .A3(_2775_),
    .ZN(_0032_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5464_ (.A1(_0002_),
    .A2(_2786_),
    .ZN(_0033_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5465_ (.A1(\title_r[12] ),
    .A2(_2574_),
    .ZN(_1866_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5466_ (.A1(\title_r[12] ),
    .A2(net152),
    .ZN(_1867_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5467_ (.A1(\title_r[9] ),
    .A2(net152),
    .Z(_1868_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5468_ (.A1(\title_r[7] ),
    .A2(net152),
    .ZN(_1869_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5469_ (.A1(\title_r[6] ),
    .A2(net156),
    .ZN(_1870_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5470_ (.A1(\title_r[6] ),
    .A2(net156),
    .ZN(_1871_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5471_ (.A1(\title_r[5] ),
    .A2(net159),
    .Z(_1872_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5472_ (.A1(\title_r[5] ),
    .A2(net159),
    .ZN(_1873_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5473_ (.A1(_1872_),
    .A2(_1873_),
    .ZN(_1874_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5474_ (.A1(\title_r[4] ),
    .A2(net161),
    .ZN(_1875_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5475_ (.A1(\title_r[3] ),
    .A2(net162),
    .ZN(_1876_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5476_ (.A1(\title_r[3] ),
    .A2(net162),
    .ZN(_1877_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5477_ (.A1(\title_r[2] ),
    .A2(\hvsync_gen.hpos[1] ),
    .ZN(_1878_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5478_ (.A1(\title_r[1] ),
    .A2(\hvsync_gen.hpos[0] ),
    .ZN(_1879_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5479_ (.A1(\title_r[1] ),
    .A2(\hvsync_gen.hpos[0] ),
    .Z(_1880_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5480_ (.A1(\title_r[0] ),
    .A2(_1880_),
    .ZN(_1881_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5481_ (.A1(_1879_),
    .A2(_1881_),
    .ZN(_1882_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5482_ (.A1(_2542_),
    .A2(_2567_),
    .ZN(_1883_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5483_ (.A1(_1878_),
    .A2(_1882_),
    .A3(_1883_),
    .ZN(_1884_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5484_ (.A1(_1878_),
    .A2(_1884_),
    .Z(_1885_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5485_ (.A1(_1877_),
    .A2(_1885_),
    .Z(_1886_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5486_ (.A1(_1876_),
    .A2(_1886_),
    .ZN(_1887_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5487_ (.A1(_2540_),
    .A2(_2569_),
    .ZN(_1888_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5488_ (.A1(_1875_),
    .A2(_1888_),
    .ZN(_1889_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5489_ (.A1(_1875_),
    .A2(_1887_),
    .A3(_1888_),
    .ZN(_1890_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5490_ (.A1(_1875_),
    .A2(_1890_),
    .ZN(_1891_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5491_ (.A1(_1874_),
    .A2(_1891_),
    .B(_1872_),
    .ZN(_1892_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5492_ (.A1(_1871_),
    .A2(_1892_),
    .B(_1870_),
    .ZN(_1893_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5493_ (.A1(_1869_),
    .A2(_1893_),
    .ZN(_1894_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5494_ (.A1(_2538_),
    .A2(net152),
    .B(_1894_),
    .ZN(_1895_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5495_ (.A1(\title_r[8] ),
    .A2(net154),
    .Z(_1896_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5496_ (.I(_1896_),
    .ZN(_1897_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5497_ (.A1(_1895_),
    .A2(_1897_),
    .ZN(_1898_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5498_ (.A1(_1868_),
    .A2(_1898_),
    .ZN(_1899_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5499_ (.A1(\title_r[11] ),
    .A2(net152),
    .Z(_1900_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5500_ (.A1(\title_r[10] ),
    .A2(_2574_),
    .ZN(_1901_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5501_ (.A1(_2535_),
    .A2(net152),
    .ZN(_1902_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5502_ (.A1(_1901_),
    .A2(_1902_),
    .ZN(_1903_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_1 _5503_ (.A1(_1868_),
    .A2(_1898_),
    .A3(_1900_),
    .A4(_1903_),
    .ZN(_1904_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5504_ (.A1(_2536_),
    .A2(_2537_),
    .B(net152),
    .ZN(_1905_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5505_ (.A1(_2534_),
    .A2(_2535_),
    .B(net152),
    .ZN(_1906_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5506_ (.A1(_1905_),
    .A2(_1906_),
    .Z(_1907_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5507_ (.A1(_1904_),
    .A2(_1907_),
    .B(_1867_),
    .ZN(_1908_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5508_ (.A1(_1866_),
    .A2(_1908_),
    .ZN(_1909_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5509_ (.A1(net63),
    .A2(_2751_),
    .ZN(_1910_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5510_ (.A1(_2565_),
    .A2(_2574_),
    .A3(_1909_),
    .ZN(_1911_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5511_ (.A1(_2755_),
    .A2(_2759_),
    .A3(_1608_),
    .ZN(_1912_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5512_ (.A1(\title_r[11] ),
    .A2(net91),
    .ZN(_1913_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5513_ (.A1(\title_r[6] ),
    .A2(net93),
    .ZN(_1914_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5514_ (.I(_1914_),
    .ZN(_1915_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5515_ (.A1(\title_r[7] ),
    .A2(net91),
    .Z(_1916_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5516_ (.A1(\title_r[5] ),
    .A2(net94),
    .ZN(_1917_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5517_ (.A1(\title_r[6] ),
    .A2(net93),
    .ZN(_1918_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5518_ (.A1(_1917_),
    .A2(_1918_),
    .ZN(_1919_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5519_ (.A1(\title_r[4] ),
    .A2(net95),
    .ZN(_1920_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5520_ (.A1(\title_r[5] ),
    .A2(net94),
    .ZN(_1921_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5521_ (.A1(_1920_),
    .A2(_1921_),
    .ZN(_1922_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5522_ (.A1(\title_r[3] ),
    .A2(net97),
    .ZN(_1923_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5523_ (.A1(\title_r[4] ),
    .A2(net95),
    .ZN(_1924_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5524_ (.A1(_1923_),
    .A2(_1924_),
    .ZN(_1925_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5525_ (.A1(\title_r[2] ),
    .A2(\hvsync_gen.vpos[1] ),
    .ZN(_1926_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5526_ (.A1(\title_r[3] ),
    .A2(net97),
    .ZN(_1927_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5527_ (.A1(_1926_),
    .A2(_1927_),
    .ZN(_1928_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5528_ (.A1(\title_r[2] ),
    .A2(\hvsync_gen.vpos[1] ),
    .ZN(_1929_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5529_ (.A1(\title_r[1] ),
    .A2(\hvsync_gen.vpos[0] ),
    .ZN(_1930_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5530_ (.A1(\title_r[1] ),
    .A2(\hvsync_gen.vpos[0] ),
    .B(\title_r[0] ),
    .ZN(_1931_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5531_ (.A1(_1930_),
    .A2(_1931_),
    .B(_1929_),
    .ZN(_1932_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5532_ (.A1(_1926_),
    .A2(_1927_),
    .Z(_1933_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5533_ (.A1(_1932_),
    .A2(_1933_),
    .B(_1928_),
    .ZN(_1934_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5534_ (.A1(_1923_),
    .A2(_1924_),
    .Z(_1935_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5535_ (.I(_1935_),
    .ZN(_1936_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5536_ (.A1(_1934_),
    .A2(_1936_),
    .ZN(_1937_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5537_ (.A1(_1925_),
    .A2(_1937_),
    .ZN(_1938_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5538_ (.A1(_1920_),
    .A2(_1921_),
    .Z(_1939_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5539_ (.I(_1939_),
    .ZN(_1940_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5540_ (.A1(_1938_),
    .A2(_1940_),
    .ZN(_1941_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5541_ (.A1(_1922_),
    .A2(_1941_),
    .ZN(_1942_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5542_ (.A1(_1917_),
    .A2(_1918_),
    .Z(_1943_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5543_ (.I(_1943_),
    .ZN(_1944_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5544_ (.A1(_1942_),
    .A2(_1944_),
    .ZN(_1945_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5545_ (.A1(_1919_),
    .A2(_1945_),
    .ZN(_1946_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5546_ (.A1(_1914_),
    .A2(_1916_),
    .ZN(_1947_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5547_ (.I(_1947_),
    .ZN(_1948_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5548_ (.A1(_1946_),
    .A2(_1948_),
    .ZN(_1949_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5549_ (.A1(_1915_),
    .A2(_1916_),
    .B(_1949_),
    .ZN(_1950_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5550_ (.A1(\title_r[10] ),
    .A2(net91),
    .ZN(_1951_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5551_ (.A1(_2534_),
    .A2(_1951_),
    .ZN(_1952_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _5552_ (.I0(\title_r[8] ),
    .I1(\title_r[7] ),
    .S(net91),
    .Z(_1953_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5553_ (.A1(\title_r[9] ),
    .A2(net91),
    .ZN(_1954_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5554_ (.A1(_2535_),
    .A2(_1954_),
    .ZN(_1955_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5555_ (.A1(_2537_),
    .A2(_2580_),
    .ZN(_1956_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5556_ (.A1(\title_r[8] ),
    .A2(net91),
    .ZN(_1957_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _5557_ (.A1(\title_r[10] ),
    .A2(\title_r[9] ),
    .A3(_1953_),
    .A4(_1956_),
    .ZN(_1958_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5558_ (.A1(\title_r[9] ),
    .A2(_1956_),
    .B(_1954_),
    .ZN(_1959_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5559_ (.A1(\title_r[8] ),
    .A2(_1954_),
    .B(_1959_),
    .ZN(_1960_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _5560_ (.I0(_2536_),
    .I1(_1955_),
    .S(_1951_),
    .Z(_1961_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5561_ (.A1(_2534_),
    .A2(_1950_),
    .A3(_1951_),
    .A4(_1958_),
    .ZN(_1962_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5562_ (.A1(\title_r[10] ),
    .A2(_1913_),
    .ZN(_1963_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5563_ (.A1(_1913_),
    .A2(_1952_),
    .B(_1963_),
    .ZN(_1964_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _5564_ (.A1(\title_r[11] ),
    .A2(net91),
    .B(_1962_),
    .C(\title_r[12] ),
    .ZN(_1965_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5565_ (.A1(\title_r[13] ),
    .A2(_1965_),
    .ZN(_1966_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai221_1 _5566_ (.A1(_2565_),
    .A2(net76),
    .B1(net46),
    .B2(_1966_),
    .C(_1912_),
    .ZN(_1967_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5567_ (.A1(_1910_),
    .A2(_1911_),
    .B(_1967_),
    .ZN(_1968_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5568_ (.A1(net167),
    .A2(_1968_),
    .ZN(_0034_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5569_ (.A1(net171),
    .A2(_1607_),
    .ZN(_1969_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5570_ (.A1(_2543_),
    .A2(net80),
    .ZN(_1970_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and4_1 _5571_ (.A1(net95),
    .A2(net97),
    .A3(net93),
    .A4(net94),
    .Z(_1971_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5572_ (.A1(net91),
    .A2(_1971_),
    .ZN(_1972_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5573_ (.A1(_2581_),
    .A2(_1972_),
    .B(\hvsync_gen.hpos[8] ),
    .ZN(_1973_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5574_ (.A1(\hvsync_gen.hpos[7] ),
    .A2(_2576_),
    .ZN(_1974_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5575_ (.A1(_2578_),
    .A2(_2758_),
    .ZN(_1975_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5576_ (.A1(net95),
    .A2(_2756_),
    .A3(_1975_),
    .ZN(_1976_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5577_ (.A1(net155),
    .A2(\title_r_pixels_in_scanline[5] ),
    .ZN(_1977_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5578_ (.A1(net162),
    .A2(\title_r_pixels_in_scanline[2] ),
    .Z(_1978_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _5579_ (.A1(\hvsync_gen.hpos[1] ),
    .A2(\title_r_pixels_in_scanline[1] ),
    .B(\title_r_pixels_in_scanline[0] ),
    .C(\hvsync_gen.hpos[0] ),
    .ZN(_1979_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5580_ (.A1(\hvsync_gen.hpos[1] ),
    .A2(\title_r_pixels_in_scanline[1] ),
    .B(_1978_),
    .ZN(_1980_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5581_ (.A1(_2570_),
    .A2(_2591_),
    .B1(_1979_),
    .B2(_1980_),
    .ZN(_1981_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5582_ (.A1(\hvsync_gen.hpos[1] ),
    .A2(\title_r_pixels_in_scanline[1] ),
    .ZN(_1982_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5583_ (.A1(\hvsync_gen.hpos[0] ),
    .A2(\title_r_pixels_in_scanline[0] ),
    .Z(_1983_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5584_ (.A1(_1978_),
    .A2(_1983_),
    .ZN(_1984_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai221_1 _5585_ (.A1(net161),
    .A2(\title_r_pixels_in_scanline[3] ),
    .B1(_1982_),
    .B2(_1984_),
    .C(_1981_),
    .ZN(_1985_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5586_ (.A1(net157),
    .A2(\title_r_pixels_in_scanline[4] ),
    .B1(\title_r_pixels_in_scanline[3] ),
    .B2(net160),
    .ZN(_1986_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5587_ (.A1(_1985_),
    .A2(_1986_),
    .ZN(_1987_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5588_ (.A1(net157),
    .A2(\title_r_pixels_in_scanline[4] ),
    .B(_1987_),
    .ZN(_1988_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5589_ (.A1(_1977_),
    .A2(_1988_),
    .ZN(_1989_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5590_ (.A1(net155),
    .A2(\title_r_pixels_in_scanline[5] ),
    .B(_1974_),
    .C(_1989_),
    .ZN(_1990_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai32_1 _5591_ (.A1(_1973_),
    .A2(_1974_),
    .A3(_1976_),
    .B1(_1990_),
    .B2(\hvsync_gen.vpos[7] ),
    .ZN(_1991_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5592_ (.A1(_2574_),
    .A2(\hvsync_gen.hpos[9] ),
    .A3(_2623_),
    .ZN(_1992_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5593_ (.A1(_2572_),
    .A2(\title_r_pixels_in_scanline[5] ),
    .ZN(_1993_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5594_ (.A1(net155),
    .A2(\title_r_pixels_in_scanline[5] ),
    .Z(_1994_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5595_ (.A1(net157),
    .A2(\title_r_pixels_in_scanline[4] ),
    .Z(_1995_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5596_ (.A1(_2568_),
    .A2(\title_r_pixels_in_scanline[0] ),
    .B(_1982_),
    .ZN(_1996_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5597_ (.A1(_2570_),
    .A2(\title_r_pixels_in_scanline[2] ),
    .B1(\title_r_pixels_in_scanline[1] ),
    .B2(_2567_),
    .ZN(_1997_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5598_ (.A1(net160),
    .A2(\title_r_pixels_in_scanline[3] ),
    .ZN(_1998_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5599_ (.A1(net162),
    .A2(_2591_),
    .B1(_1996_),
    .B2(_1997_),
    .ZN(_1999_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5600_ (.A1(_2569_),
    .A2(\title_r_pixels_in_scanline[3] ),
    .B1(_1998_),
    .B2(_1999_),
    .ZN(_2000_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5601_ (.A1(_1995_),
    .A2(_2000_),
    .ZN(_2001_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5602_ (.A1(_2571_),
    .A2(\title_r_pixels_in_scanline[4] ),
    .B(_2001_),
    .ZN(_2002_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5603_ (.A1(_1994_),
    .A2(_2002_),
    .B(_1993_),
    .ZN(_2003_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5604_ (.A1(_1978_),
    .A2(_1983_),
    .ZN(_2004_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5605_ (.A1(_1994_),
    .A2(_1995_),
    .ZN(_2005_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5606_ (.A1(_1982_),
    .A2(_1998_),
    .A3(_2004_),
    .A4(_2005_),
    .ZN(_2006_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _5607_ (.A1(\hvsync_gen.hpos[8] ),
    .A2(_2580_),
    .B(\hvsync_gen.hpos[7] ),
    .C(\hvsync_gen.hpos[9] ),
    .ZN(_2007_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_1 _5608_ (.A1(net153),
    .A2(\hvsync_gen.vpos[7] ),
    .A3(_2623_),
    .A4(_2007_),
    .ZN(_2008_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5609_ (.A1(_2003_),
    .A2(_2008_),
    .Z(_2009_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5610_ (.A1(_1991_),
    .A2(_1992_),
    .B1(_2006_),
    .B2(_2009_),
    .ZN(_2010_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5611_ (.A1(\ppp_y[4] ),
    .A2(\ppp_y[5] ),
    .ZN(_2011_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5612_ (.A1(\ppp_y[4] ),
    .A2(\ppp_y[3] ),
    .A3(\ppp_y[5] ),
    .ZN(_2012_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5613_ (.I(_2012_),
    .ZN(_2013_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5614_ (.A1(_2010_),
    .A2(_2012_),
    .ZN(_2014_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _5615_ (.A1(_2543_),
    .A2(net80),
    .A3(_2014_),
    .ZN(_2015_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5616_ (.A1(\ppp_y[7] ),
    .A2(\ppp_y[6] ),
    .ZN(_2016_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5617_ (.A1(_2779_),
    .A2(_2010_),
    .Z(_2017_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5618_ (.A1(_2016_),
    .A2(_2017_),
    .Z(_2018_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5619_ (.A1(_2543_),
    .A2(net71),
    .ZN(_2019_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5620_ (.A1(net111),
    .A2(_0224_),
    .B(\ppp_y[7] ),
    .ZN(_2020_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _5621_ (.A1(_2543_),
    .A2(_2594_),
    .A3(net71),
    .A4(_2011_),
    .ZN(_2021_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5622_ (.A1(_2633_),
    .A2(_2021_),
    .ZN(_2022_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _5623_ (.A1(_2018_),
    .A2(_2019_),
    .A3(_2020_),
    .B(_2022_),
    .ZN(_2023_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5624_ (.A1(\ppp_y[3] ),
    .A2(\ppp_y[1] ),
    .A3(\ppp_y[2] ),
    .ZN(_2024_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5625_ (.A1(_2011_),
    .A2(_2024_),
    .B(_2634_),
    .ZN(_2025_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5626_ (.A1(\frame_counter[9] ),
    .A2(_0225_),
    .ZN(_2026_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5627_ (.A1(_2543_),
    .A2(_0224_),
    .ZN(_2027_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5628_ (.A1(_2016_),
    .A2(_2026_),
    .ZN(_2028_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5629_ (.A1(_1970_),
    .A2(_2023_),
    .A3(_2025_),
    .A4(_2028_),
    .ZN(_2029_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5630_ (.A1(_2015_),
    .A2(_2029_),
    .B(_1969_),
    .ZN(_0035_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _5631_ (.A1(net111),
    .A2(_0224_),
    .A3(_2017_),
    .Z(_2030_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5632_ (.A1(_2020_),
    .A2(_2030_),
    .B(_2638_),
    .ZN(_2031_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5633_ (.A1(_2633_),
    .A2(_2019_),
    .ZN(_2032_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5634_ (.A1(\ppp_y[6] ),
    .A2(_2638_),
    .B(_2031_),
    .C(_2032_),
    .ZN(_2033_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5635_ (.A1(_2594_),
    .A2(_2011_),
    .A3(_2024_),
    .ZN(_2034_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5636_ (.A1(\ppp_y[0] ),
    .A2(_2634_),
    .A3(_2034_),
    .ZN(_2035_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5637_ (.A1(_2033_),
    .A2(_2035_),
    .ZN(_2036_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5638_ (.A1(_1970_),
    .A2(_2036_),
    .ZN(_2037_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5639_ (.A1(_2015_),
    .A2(_2037_),
    .B(_1969_),
    .ZN(_0036_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _5640_ (.I0(net102),
    .I1(\ppp_y[5] ),
    .S(_2016_),
    .Z(_2038_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5641_ (.I(_2038_),
    .ZN(_2039_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5642_ (.A1(\ppp_x[6] ),
    .A2(_2020_),
    .B1(_2030_),
    .B2(_2039_),
    .ZN(_2040_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5643_ (.A1(_2636_),
    .A2(_2040_),
    .ZN(_2041_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _5644_ (.A1(\ppp_y[4] ),
    .A2(\ppp_y[3] ),
    .A3(\dot[7] ),
    .A4(_2021_),
    .ZN(_2042_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5645_ (.A1(\ppp_y[5] ),
    .A2(_2637_),
    .ZN(_2043_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _5646_ (.A1(_2027_),
    .A2(_2041_),
    .A3(_2042_),
    .A4(_2043_),
    .ZN(_2044_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5647_ (.A1(net111),
    .A2(\frame_counter[8] ),
    .B1(_2027_),
    .B2(_2038_),
    .C(_2044_),
    .ZN(_2045_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5648_ (.A1(_2015_),
    .A2(_2045_),
    .B(_1969_),
    .ZN(_0037_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5649_ (.A1(net111),
    .A2(_0224_),
    .B(\ppp_y[6] ),
    .ZN(_2046_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5650_ (.A1(_2021_),
    .A2(_2026_),
    .ZN(_2047_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _5651_ (.A1(_2018_),
    .A2(_2019_),
    .A3(_2046_),
    .B(_2047_),
    .ZN(_2048_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _5652_ (.A1(_2635_),
    .A2(_1970_),
    .A3(_2028_),
    .A4(_2048_),
    .ZN(_2049_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _5653_ (.A1(\ppp_y[0] ),
    .A2(\ppp_y[2] ),
    .A3(_2634_),
    .A4(_2013_),
    .ZN(_2050_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5654_ (.A1(_2049_),
    .A2(_2050_),
    .Z(_2051_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5655_ (.A1(_2015_),
    .A2(_2051_),
    .B(_1969_),
    .ZN(_0038_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _5656_ (.A1(_2637_),
    .A2(_2030_),
    .A3(_2046_),
    .B(_2043_),
    .ZN(_2052_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5657_ (.A1(_2032_),
    .A2(_2052_),
    .ZN(_2053_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5658_ (.A1(_2035_),
    .A2(_2053_),
    .ZN(_2054_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5659_ (.A1(_1970_),
    .A2(_2054_),
    .ZN(_2055_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5660_ (.A1(_2015_),
    .A2(_2055_),
    .B(_1969_),
    .ZN(_0039_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _5661_ (.I0(\dot[5] ),
    .I1(\ppp_y[4] ),
    .S(_2016_),
    .Z(_2056_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5662_ (.I(_2056_),
    .ZN(_2057_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5663_ (.A1(\ppp_x[5] ),
    .A2(_2046_),
    .B1(_2057_),
    .B2(_2030_),
    .ZN(_2058_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5664_ (.A1(\ppp_y[4] ),
    .A2(_2637_),
    .B1(_2058_),
    .B2(_2636_),
    .C(_2026_),
    .ZN(_2059_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5665_ (.A1(_2026_),
    .A2(_2057_),
    .B(_2059_),
    .ZN(_2060_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5666_ (.A1(_2635_),
    .A2(_1970_),
    .A3(_2060_),
    .ZN(_2061_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5667_ (.A1(_2015_),
    .A2(_2061_),
    .B(_1969_),
    .ZN(_0040_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5668_ (.A1(\r1[8] ),
    .A2(\r1[9] ),
    .A3(_2952_),
    .ZN(_2062_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5669_ (.A1(\r1[12] ),
    .A2(\r1[13] ),
    .Z(_2063_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5670_ (.A1(net98),
    .A2(\r1[11] ),
    .A3(_2063_),
    .ZN(_2064_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5671_ (.A1(\r1[2] ),
    .A2(\r1[3] ),
    .ZN(_2065_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5672_ (.A1(_2062_),
    .A2(_2064_),
    .A3(_2065_),
    .ZN(_2066_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5673_ (.A1(\r1[4] ),
    .A2(\r1[5] ),
    .Z(_2067_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5674_ (.A1(_2614_),
    .A2(\r1[7] ),
    .A3(_2067_),
    .ZN(_2068_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5675_ (.A1(_2618_),
    .A2(\r1[17] ),
    .ZN(_2069_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5676_ (.A1(\r1[16] ),
    .A2(\r1[17] ),
    .ZN(_2070_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5677_ (.A1(_2609_),
    .A2(\r1[1] ),
    .A3(_2070_),
    .ZN(_2071_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5678_ (.A1(_2066_),
    .A2(_2068_),
    .A3(_2071_),
    .ZN(_2072_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5679_ (.A1(\noise_counter[2] ),
    .A2(\noise_counter[1] ),
    .ZN(_2073_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5680_ (.A1(net58),
    .A2(_2072_),
    .A3(_2073_),
    .ZN(_2074_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5681_ (.A1(noise),
    .A2(_2074_),
    .Z(_2075_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5682_ (.A1(net169),
    .A2(_2075_),
    .Z(_0041_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _5683_ (.A1(\noise_counter[2] ),
    .A2(\noise_counter[1] ),
    .A3(\noise_counter[0] ),
    .B(net59),
    .ZN(_2076_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5684_ (.A1(\noise_counter[0] ),
    .A2(net59),
    .B(_2076_),
    .C(net169),
    .ZN(_2077_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5685_ (.I(_2077_),
    .ZN(_0042_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5686_ (.A1(\noise_counter[1] ),
    .A2(net59),
    .ZN(_2078_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5687_ (.A1(\noise_counter[0] ),
    .A2(_2073_),
    .ZN(_2079_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _5688_ (.A1(net59),
    .A2(_2079_),
    .B(_2078_),
    .C(net164),
    .ZN(_0043_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _5689_ (.A1(\noise_counter[2] ),
    .A2(net169),
    .A3(net58),
    .Z(_0044_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5690_ (.A1(_2563_),
    .A2(\note2_freq[1] ),
    .B1(\note2_freq[0] ),
    .B2(_2564_),
    .ZN(_2080_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5691_ (.A1(_2562_),
    .A2(\note2_freq[3] ),
    .B1(\note2_freq[1] ),
    .B2(_2563_),
    .ZN(_2081_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5692_ (.A1(\note2_counter[2] ),
    .A2(_2080_),
    .A3(_2081_),
    .ZN(_2082_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5693_ (.A1(_2562_),
    .A2(\note2_freq[3] ),
    .Z(_2083_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5694_ (.A1(_2561_),
    .A2(\note2_freq[4] ),
    .B1(_2082_),
    .B2(_2083_),
    .ZN(_2084_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5695_ (.A1(_2560_),
    .A2(\note2_freq[5] ),
    .B1(\note2_freq[4] ),
    .B2(_2561_),
    .ZN(_2085_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5696_ (.A1(_2559_),
    .A2(\note2_freq[6] ),
    .B1(\note2_freq[5] ),
    .B2(_2560_),
    .ZN(_2086_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5697_ (.A1(_2084_),
    .A2(_2085_),
    .B(_2086_),
    .ZN(_2087_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _5698_ (.A1(_2558_),
    .A2(\note2_freq[7] ),
    .B1(\note2_freq[6] ),
    .B2(_2559_),
    .C(_2087_),
    .ZN(_2088_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5699_ (.A1(_2557_),
    .A2(\note2_freq[8] ),
    .B1(\note2_freq[7] ),
    .B2(_2558_),
    .ZN(_2089_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5700_ (.A1(\note2_counter[8] ),
    .A2(_2585_),
    .B1(_2088_),
    .B2(_2089_),
    .ZN(_2090_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5701_ (.A1(net58),
    .A2(_2090_),
    .Z(_2091_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5702_ (.A1(net169),
    .A2(_2091_),
    .ZN(_2092_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5703_ (.A1(\note2_counter[0] ),
    .A2(net59),
    .ZN(_2093_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5704_ (.A1(_2092_),
    .A2(_2093_),
    .ZN(_0045_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5705_ (.A1(\note2_counter[0] ),
    .A2(net59),
    .B(\note2_counter[1] ),
    .ZN(_2094_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _5706_ (.A1(_2563_),
    .A2(_2564_),
    .A3(net58),
    .ZN(_2095_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5707_ (.A1(_2092_),
    .A2(_2094_),
    .A3(_2095_),
    .ZN(_0046_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5708_ (.A1(\note2_counter[2] ),
    .A2(_2095_),
    .ZN(_2096_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5709_ (.A1(_2092_),
    .A2(_2096_),
    .ZN(_0047_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5710_ (.A1(\note2_counter[2] ),
    .A2(_2095_),
    .B(\note2_counter[3] ),
    .ZN(_2097_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and4_1 _5711_ (.A1(\note2_counter[3] ),
    .A2(\note2_counter[2] ),
    .A3(\note2_counter[1] ),
    .A4(\note2_counter[0] ),
    .Z(_2098_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5712_ (.A1(net59),
    .A2(_2098_),
    .Z(_2099_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5713_ (.A1(_2092_),
    .A2(_2097_),
    .A3(_2099_),
    .ZN(_0048_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5714_ (.A1(\note2_counter[4] ),
    .A2(_2099_),
    .ZN(_2100_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5715_ (.A1(\note2_counter[4] ),
    .A2(_2099_),
    .Z(_2101_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5716_ (.A1(_2092_),
    .A2(_2100_),
    .A3(_2101_),
    .ZN(_0049_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _5717_ (.A1(\note2_counter[5] ),
    .A2(\note2_counter[4] ),
    .A3(_2098_),
    .Z(_2102_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5718_ (.A1(\note2_counter[5] ),
    .A2(\note2_counter[4] ),
    .A3(_2098_),
    .ZN(_2103_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5719_ (.A1(\note2_counter[5] ),
    .A2(net58),
    .B1(_2090_),
    .B2(_2103_),
    .ZN(_2104_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5720_ (.A1(\note2_counter[5] ),
    .A2(_2101_),
    .B(net170),
    .ZN(_2105_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5721_ (.A1(_2104_),
    .A2(_2105_),
    .ZN(_0050_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5722_ (.A1(_2559_),
    .A2(net58),
    .A3(_2103_),
    .ZN(_2106_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5723_ (.A1(net59),
    .A2(_2102_),
    .B(\note2_counter[6] ),
    .ZN(_2107_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5724_ (.A1(_2092_),
    .A2(_2106_),
    .A3(_2107_),
    .ZN(_0051_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5725_ (.A1(\note2_counter[7] ),
    .A2(\note2_counter[6] ),
    .A3(_2102_),
    .ZN(_2108_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5726_ (.A1(\note2_counter[7] ),
    .A2(net58),
    .B1(_2090_),
    .B2(_2108_),
    .ZN(_2109_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5727_ (.A1(\note2_counter[7] ),
    .A2(_2106_),
    .B(net170),
    .ZN(_2110_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5728_ (.A1(_2109_),
    .A2(_2110_),
    .ZN(_0052_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5729_ (.A1(\note2_counter[7] ),
    .A2(_2106_),
    .ZN(_2111_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5730_ (.A1(_2557_),
    .A2(_2111_),
    .ZN(_2112_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5731_ (.A1(_2092_),
    .A2(_2112_),
    .ZN(_0053_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5732_ (.A1(note2),
    .A2(_2091_),
    .Z(_2113_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5733_ (.A1(net164),
    .A2(_2113_),
    .ZN(_0054_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5734_ (.A1(\note_counter[6] ),
    .A2(_2586_),
    .ZN(_2114_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5735_ (.A1(\note_counter[5] ),
    .A2(_2587_),
    .B1(_2588_),
    .B2(\note_counter[4] ),
    .ZN(_2115_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5736_ (.A1(_2555_),
    .A2(\note_freq[2] ),
    .ZN(_2116_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5737_ (.A1(\note_counter[1] ),
    .A2(_2116_),
    .B(\note_counter[3] ),
    .ZN(_2117_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5738_ (.A1(_2556_),
    .A2(\note_freq[0] ),
    .ZN(_2118_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5739_ (.A1(_2554_),
    .A2(\note_freq[7] ),
    .ZN(_2119_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5740_ (.A1(_2556_),
    .A2(\note_freq[0] ),
    .B(_2119_),
    .ZN(_2120_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5741_ (.A1(\note_counter[1] ),
    .A2(_2589_),
    .B1(_2118_),
    .B2(_2120_),
    .C(_2116_),
    .ZN(_2121_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5742_ (.A1(_2555_),
    .A2(\note_freq[2] ),
    .B1(_2117_),
    .B2(\note_freq[1] ),
    .C(_2121_),
    .ZN(_2122_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5743_ (.A1(\note_counter[4] ),
    .A2(_2588_),
    .B1(_2589_),
    .B2(\note_counter[3] ),
    .C(_2122_),
    .ZN(_2123_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5744_ (.A1(_2115_),
    .A2(_2123_),
    .ZN(_2124_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5745_ (.A1(\note_counter[6] ),
    .A2(_2586_),
    .B1(_2587_),
    .B2(\note_counter[5] ),
    .C(_2124_),
    .ZN(_2125_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5746_ (.A1(_2554_),
    .A2(\note_freq[7] ),
    .B1(_2114_),
    .B2(_2125_),
    .ZN(_2126_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _5747_ (.A1(_2753_),
    .A2(_2119_),
    .A3(_2126_),
    .ZN(_2127_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _5748_ (.A1(net170),
    .A2(_2127_),
    .ZN(_2128_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5749_ (.A1(\note_counter[0] ),
    .A2(_2753_),
    .ZN(_2129_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5750_ (.A1(_2128_),
    .A2(_2129_),
    .ZN(_0055_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _5751_ (.A1(\note_counter[1] ),
    .A2(\note_counter[0] ),
    .A3(_2753_),
    .Z(_2130_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5752_ (.A1(\note_counter[0] ),
    .A2(_2753_),
    .B(\note_counter[1] ),
    .ZN(_2131_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5753_ (.A1(_2128_),
    .A2(_2130_),
    .A3(_2131_),
    .ZN(_0056_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5754_ (.A1(\note_counter[2] ),
    .A2(_2130_),
    .Z(_2132_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5755_ (.A1(\note_counter[2] ),
    .A2(_2130_),
    .ZN(_2133_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5756_ (.A1(_2128_),
    .A2(_2132_),
    .A3(_2133_),
    .ZN(_0057_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5757_ (.A1(\note_counter[3] ),
    .A2(_2132_),
    .Z(_2134_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5758_ (.A1(\note_counter[3] ),
    .A2(_2132_),
    .ZN(_2135_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5759_ (.A1(_2128_),
    .A2(_2134_),
    .A3(_2135_),
    .ZN(_0058_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5760_ (.A1(\note_counter[4] ),
    .A2(_2134_),
    .Z(_2136_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5761_ (.A1(\note_counter[4] ),
    .A2(_2134_),
    .ZN(_2137_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5762_ (.A1(_2128_),
    .A2(_2136_),
    .A3(_2137_),
    .ZN(_0059_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5763_ (.A1(\note_counter[5] ),
    .A2(_2136_),
    .Z(_2138_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5764_ (.A1(\note_counter[5] ),
    .A2(_2136_),
    .ZN(_2139_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5765_ (.A1(_2128_),
    .A2(_2138_),
    .A3(_2139_),
    .ZN(_0060_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5766_ (.A1(\note_counter[6] ),
    .A2(_2138_),
    .ZN(_2140_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5767_ (.A1(\note_counter[6] ),
    .A2(_2138_),
    .ZN(_2141_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5768_ (.A1(_2128_),
    .A2(_2141_),
    .ZN(_0061_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5769_ (.A1(_2554_),
    .A2(_2140_),
    .ZN(_2142_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5770_ (.A1(_2128_),
    .A2(_2142_),
    .ZN(_0062_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5771_ (.A1(_2553_),
    .A2(_2127_),
    .B(net170),
    .ZN(_2143_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5772_ (.A1(_2553_),
    .A2(_2127_),
    .B(_2143_),
    .ZN(_0063_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5773_ (.A1(_2567_),
    .A2(_2568_),
    .ZN(_2144_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _5774_ (.A1(_2567_),
    .A2(_2568_),
    .A3(_2569_),
    .A4(_2570_),
    .ZN(_2145_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5775_ (.A1(net157),
    .A2(_2145_),
    .Z(_2146_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5776_ (.A1(\hvsync_gen.hpos[9] ),
    .A2(_2629_),
    .A3(_1974_),
    .A4(_2146_),
    .ZN(_2147_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_1 _5777_ (.I(_2147_),
    .ZN(_2148_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5778_ (.A1(net167),
    .A2(_2148_),
    .ZN(_2149_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5779_ (.A1(net171),
    .A2(_2147_),
    .ZN(_2150_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5780_ (.A1(\hvsync_gen.hpos[0] ),
    .A2(net27),
    .ZN(_0064_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5781_ (.A1(_2748_),
    .A2(_2144_),
    .A3(net27),
    .ZN(_0065_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5782_ (.A1(net162),
    .A2(_2144_),
    .B(net171),
    .ZN(_2151_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5783_ (.A1(net162),
    .A2(_2144_),
    .B(_2151_),
    .ZN(_0066_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5784_ (.A1(net162),
    .A2(_2144_),
    .B(net160),
    .ZN(_2152_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5785_ (.A1(net167),
    .A2(_2145_),
    .A3(_2152_),
    .ZN(_0067_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5786_ (.A1(net157),
    .A2(_2145_),
    .B(net171),
    .ZN(_2153_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5787_ (.A1(_2146_),
    .A2(_2153_),
    .ZN(_0068_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5788_ (.A1(net155),
    .A2(_2146_),
    .Z(_2154_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5789_ (.A1(net155),
    .A2(_2146_),
    .ZN(_2155_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5790_ (.A1(_2150_),
    .A2(_2154_),
    .A3(_2155_),
    .ZN(_0069_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5791_ (.A1(net153),
    .A2(_2154_),
    .ZN(_2156_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5792_ (.A1(net153),
    .A2(_2154_),
    .Z(_2157_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5793_ (.A1(net27),
    .A2(_2156_),
    .A3(_2157_),
    .ZN(_0070_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5794_ (.A1(\hvsync_gen.hpos[7] ),
    .A2(_2157_),
    .ZN(_2158_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5795_ (.A1(_2628_),
    .A2(_2145_),
    .Z(_2159_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5796_ (.A1(net27),
    .A2(_2158_),
    .A3(_2159_),
    .ZN(_0071_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5797_ (.A1(\hvsync_gen.hpos[8] ),
    .A2(_2159_),
    .ZN(_2160_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5798_ (.A1(\hvsync_gen.hpos[8] ),
    .A2(_2159_),
    .ZN(_2161_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5799_ (.A1(net27),
    .A2(_2161_),
    .ZN(_0072_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5800_ (.A1(_2575_),
    .A2(_2160_),
    .ZN(_2162_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5801_ (.A1(_2150_),
    .A2(_2162_),
    .ZN(_0073_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5802_ (.A1(net167),
    .A2(net82),
    .ZN(_0074_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5803_ (.A1(net171),
    .A2(hsync),
    .Z(_0075_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5804_ (.A1(net144),
    .A2(_2762_),
    .B(net170),
    .ZN(_2163_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5805_ (.A1(_2763_),
    .A2(_2163_),
    .ZN(_0076_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5806_ (.A1(net136),
    .A2(_2763_),
    .B(net172),
    .ZN(_2164_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5807_ (.A1(_2764_),
    .A2(_2164_),
    .ZN(_0077_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5808_ (.A1(net131),
    .A2(_2764_),
    .ZN(_2165_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5809_ (.A1(net166),
    .A2(_2766_),
    .A3(_2165_),
    .ZN(_0078_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5810_ (.A1(_2545_),
    .A2(_2781_),
    .B(_2544_),
    .ZN(_2166_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _5811_ (.A1(\frame_counter[8] ),
    .A2(\frame_counter[7] ),
    .A3(net112),
    .A4(_2771_),
    .ZN(_2167_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5812_ (.A1(net172),
    .A2(_2166_),
    .A3(_2167_),
    .ZN(_2168_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5813_ (.I(_2168_),
    .ZN(_0084_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5814_ (.A1(_2543_),
    .A2(_2167_),
    .ZN(_2169_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5815_ (.A1(net168),
    .A2(_2169_),
    .ZN(_0085_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5816_ (.A1(frame_counter_frac),
    .A2(_2761_),
    .B(net171),
    .ZN(_2170_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5817_ (.A1(_2762_),
    .A2(_2170_),
    .ZN(_0086_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5818_ (.A1(frame_counter_frac),
    .A2(net163),
    .B(net160),
    .ZN(_2171_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5819_ (.A1(net143),
    .A2(net160),
    .B1(net157),
    .B2(net137),
    .ZN(_2172_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _5820_ (.A1(net143),
    .A2(net160),
    .B(net163),
    .C(frame_counter_frac),
    .ZN(_2173_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5821_ (.A1(net137),
    .A2(net157),
    .B1(net156),
    .B2(net130),
    .ZN(_2174_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5822_ (.A1(_2172_),
    .A2(_2173_),
    .B(_2174_),
    .ZN(_2175_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai221_1 _5823_ (.A1(net130),
    .A2(net155),
    .B1(net153),
    .B2(net127),
    .C(_2175_),
    .ZN(_2176_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _5824_ (.A1(net126),
    .A2(net154),
    .B(\hvsync_gen.vpos[9] ),
    .C(_2747_),
    .ZN(_2177_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _5825_ (.A1(_2566_),
    .A2(_2577_),
    .ZN(_2178_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5826_ (.A1(net97),
    .A2(_2178_),
    .B(net95),
    .ZN(_2179_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _5827_ (.A1(\hvsync_gen.vpos[1] ),
    .A2(net97),
    .B(_2756_),
    .C(net95),
    .ZN(_2180_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5828_ (.A1(_2582_),
    .A2(_2180_),
    .B(_2177_),
    .C(_2176_),
    .ZN(_2181_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5829_ (.A1(net130),
    .A2(\hvsync_gen.hpos[7] ),
    .ZN(_2182_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5830_ (.A1(net160),
    .A2(net157),
    .B(frame_counter_frac),
    .ZN(_2183_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5831_ (.A1(net160),
    .A2(net157),
    .B1(net156),
    .B2(net143),
    .ZN(_2184_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5832_ (.A1(net143),
    .A2(net156),
    .ZN(_2185_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5833_ (.A1(_2551_),
    .A2(_2574_),
    .B1(_2183_),
    .B2(_2184_),
    .C(_2185_),
    .ZN(_2186_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5834_ (.A1(net130),
    .A2(\hvsync_gen.hpos[7] ),
    .B1(net153),
    .B2(net142),
    .C(_2186_),
    .ZN(_2187_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5835_ (.A1(note),
    .A2(_2575_),
    .A3(\hvsync_gen.hpos[8] ),
    .ZN(_2188_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5836_ (.A1(\frame_counter[9] ),
    .A2(_0224_),
    .B1(_2182_),
    .B2(_2187_),
    .ZN(_2189_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5837_ (.A1(_2629_),
    .A2(_0203_),
    .ZN(_2190_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5838_ (.A1(note2),
    .A2(\hvsync_gen.hpos[9] ),
    .ZN(_2191_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5839_ (.A1(frame_counter_frac),
    .A2(net163),
    .B1(net158),
    .B2(net143),
    .ZN(_2192_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5840_ (.A1(_2171_),
    .A2(_2192_),
    .ZN(_2193_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5841_ (.A1(net143),
    .A2(net158),
    .B(_2193_),
    .ZN(_2194_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5842_ (.A1(_2551_),
    .A2(_2572_),
    .B(_2194_),
    .ZN(_2195_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai221_1 _5843_ (.A1(net142),
    .A2(net155),
    .B1(net153),
    .B2(net130),
    .C(_2195_),
    .ZN(_2196_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5844_ (.A1(noise),
    .A2(_2625_),
    .ZN(_2197_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _5845_ (.A1(net130),
    .A2(net153),
    .B(\hvsync_gen.hpos[9] ),
    .C(_2197_),
    .ZN(_2198_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _5846_ (.A1(_0202_),
    .A2(_1970_),
    .A3(_2196_),
    .A4(_2198_),
    .ZN(_2199_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _5847_ (.A1(_2746_),
    .A2(_2190_),
    .A3(_2191_),
    .B(_2199_),
    .ZN(_2200_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5848_ (.I(_2200_),
    .ZN(_2201_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5849_ (.A1(_2188_),
    .A2(_2189_),
    .B(_2201_),
    .C(_2181_),
    .ZN(_2202_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5850_ (.A1(net171),
    .A2(_2202_),
    .Z(_0087_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5851_ (.A1(net112),
    .A2(\hvsync_gen.hpos[7] ),
    .B(net154),
    .ZN(_2203_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5852_ (.A1(_2879_),
    .A2(_2203_),
    .ZN(_2204_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5853_ (.A1(net142),
    .A2(_2567_),
    .B1(_2568_),
    .B2(net143),
    .ZN(_2205_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5854_ (.A1(_2551_),
    .A2(\hvsync_gen.hpos[1] ),
    .B1(net163),
    .B2(_2550_),
    .C(_2205_),
    .ZN(_2206_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5855_ (.A1(net126),
    .A2(_2569_),
    .B1(_2570_),
    .B2(net130),
    .C(_2206_),
    .ZN(_2207_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5856_ (.A1(_2549_),
    .A2(net161),
    .B1(net158),
    .B2(net122),
    .C(_2207_),
    .ZN(_2208_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5857_ (.A1(net122),
    .A2(net158),
    .B1(net156),
    .B2(net57),
    .ZN(_2209_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai222_1 _5858_ (.A1(_2572_),
    .A2(net56),
    .B1(_2208_),
    .B2(_2209_),
    .C1(_2879_),
    .C2(_2574_),
    .ZN(_2210_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5859_ (.A1(_2204_),
    .A2(_2210_),
    .ZN(_2211_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5860_ (.A1(\hvsync_gen.hpos[7] ),
    .A2(_2876_),
    .B(\hvsync_gen.hpos[8] ),
    .ZN(_2212_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _5861_ (.A1(_2576_),
    .A2(_2877_),
    .B1(_2211_),
    .B2(_2212_),
    .ZN(_2213_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _5862_ (.A1(\hvsync_gen.hpos[9] ),
    .A2(_2213_),
    .ZN(_2214_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _5863_ (.A1(\hvsync_gen.hpos[9] ),
    .A2(_2213_),
    .Z(_2215_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5864_ (.A1(net144),
    .A2(\r1[0] ),
    .ZN(_2216_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5865_ (.A1(net144),
    .A2(\r1[0] ),
    .Z(_2217_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5866_ (.A1(net84),
    .A2(\r1[0] ),
    .A3(net13),
    .ZN(_2218_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5867_ (.A1(_2214_),
    .A2(_2217_),
    .B(net34),
    .ZN(_2219_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5868_ (.A1(net90),
    .A2(_2609_),
    .A3(net28),
    .ZN(_2220_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5869_ (.A1(_2609_),
    .A2(net28),
    .B(_2220_),
    .ZN(_2221_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5870_ (.A1(_2218_),
    .A2(_2219_),
    .B1(_2221_),
    .B2(net34),
    .C(net166),
    .ZN(_0088_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5871_ (.A1(_2610_),
    .A2(_0230_),
    .ZN(_2222_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5872_ (.A1(\r1[0] ),
    .A2(_2222_),
    .ZN(_2223_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5873_ (.A1(\r1[0] ),
    .A2(_2222_),
    .Z(_2224_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5874_ (.A1(net28),
    .A2(_2223_),
    .A3(_2224_),
    .ZN(_2225_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _5875_ (.A1(net89),
    .A2(net28),
    .ZN(_2226_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5876_ (.A1(\r1[1] ),
    .A2(_2226_),
    .B(net39),
    .ZN(_2227_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5877_ (.A1(net84),
    .A2(\r1[1] ),
    .A3(net13),
    .ZN(_2228_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5878_ (.A1(net137),
    .A2(\r1[1] ),
    .ZN(_2229_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5879_ (.A1(net137),
    .A2(\r1[1] ),
    .ZN(_2230_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5880_ (.A1(_2551_),
    .A2(_2610_),
    .A3(_2216_),
    .ZN(_2231_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5881_ (.A1(_2214_),
    .A2(_2231_),
    .B(net34),
    .ZN(_2232_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5882_ (.A1(_2225_),
    .A2(_2227_),
    .B1(_2228_),
    .B2(_2232_),
    .C(net166),
    .ZN(_0089_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5883_ (.A1(_2611_),
    .A2(net19),
    .ZN(_2233_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5884_ (.A1(_2611_),
    .A2(net19),
    .ZN(_2234_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5885_ (.A1(_2610_),
    .A2(_0231_),
    .B(_2223_),
    .ZN(_2235_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5886_ (.A1(\r1[2] ),
    .A2(net19),
    .A3(_2235_),
    .ZN(_2236_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5887_ (.A1(net84),
    .A2(\r1[2] ),
    .ZN(_2237_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5888_ (.A1(net45),
    .A2(_2237_),
    .B(net38),
    .ZN(_2238_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5889_ (.A1(net45),
    .A2(_2236_),
    .B(_2238_),
    .ZN(_2239_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5890_ (.A1(net131),
    .A2(\r1[2] ),
    .Z(_2240_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5891_ (.A1(_2216_),
    .A2(_2230_),
    .B(_2229_),
    .ZN(_2241_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5892_ (.A1(_2240_),
    .A2(_2241_),
    .ZN(_2242_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5893_ (.A1(_2240_),
    .A2(_2241_),
    .ZN(_2243_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5894_ (.A1(_2214_),
    .A2(_2243_),
    .ZN(_2244_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5895_ (.A1(net13),
    .A2(_2237_),
    .ZN(_2245_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5896_ (.A1(net39),
    .A2(_2244_),
    .A3(_2245_),
    .ZN(_2246_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5897_ (.A1(_2239_),
    .A2(_2246_),
    .B(net166),
    .ZN(_0090_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5898_ (.A1(_2234_),
    .A2(_2235_),
    .B(_2233_),
    .ZN(_2247_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5899_ (.A1(\r1[3] ),
    .A2(net18),
    .ZN(_2248_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5900_ (.A1(\r1[3] ),
    .A2(net18),
    .ZN(_2249_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5901_ (.A1(\r1[3] ),
    .A2(net18),
    .A3(_2247_),
    .ZN(_2250_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5902_ (.A1(net90),
    .A2(_2612_),
    .B(net45),
    .ZN(_2251_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5903_ (.A1(net45),
    .A2(_2250_),
    .B(_2251_),
    .C(net34),
    .ZN(_2252_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5904_ (.A1(net127),
    .A2(\r1[3] ),
    .Z(_2253_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5905_ (.A1(_2550_),
    .A2(_2611_),
    .B(_2242_),
    .ZN(_2254_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5906_ (.A1(_2253_),
    .A2(_2254_),
    .ZN(_2255_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5907_ (.A1(_2253_),
    .A2(_2254_),
    .Z(_2256_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5908_ (.A1(net90),
    .A2(_2612_),
    .B(net13),
    .ZN(_2257_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5909_ (.A1(net13),
    .A2(_2256_),
    .B(_2257_),
    .C(net38),
    .ZN(_2258_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5910_ (.A1(_2252_),
    .A2(_2258_),
    .B(net166),
    .ZN(_0091_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5911_ (.A1(net122),
    .A2(_2613_),
    .ZN(_2259_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5912_ (.A1(_2548_),
    .A2(\r1[4] ),
    .ZN(_2260_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5913_ (.A1(_2259_),
    .A2(_2260_),
    .ZN(_2261_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5914_ (.A1(_2549_),
    .A2(_2612_),
    .B(_2255_),
    .ZN(_2262_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5915_ (.A1(_2261_),
    .A2(_2262_),
    .ZN(_2263_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5916_ (.A1(_2214_),
    .A2(_2263_),
    .ZN(_2264_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5917_ (.A1(net90),
    .A2(_2613_),
    .ZN(_2265_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5918_ (.A1(_2214_),
    .A2(_2265_),
    .B(_2264_),
    .C(net38),
    .ZN(_2266_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5919_ (.A1(_2247_),
    .A2(_2249_),
    .B(_2248_),
    .ZN(_2267_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5920_ (.A1(_2613_),
    .A2(_0330_),
    .ZN(_2268_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5921_ (.A1(_2613_),
    .A2(_0330_),
    .ZN(_2269_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5922_ (.A1(_2613_),
    .A2(_0330_),
    .A3(_2267_),
    .ZN(_2270_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5923_ (.A1(net29),
    .A2(_2270_),
    .ZN(_2271_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5924_ (.A1(net29),
    .A2(_2265_),
    .B(_2271_),
    .C(net34),
    .ZN(_2272_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5925_ (.A1(_2266_),
    .A2(_2272_),
    .B(net168),
    .ZN(_0092_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5926_ (.A1(net84),
    .A2(\r1[5] ),
    .ZN(_2273_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5927_ (.A1(net45),
    .A2(_2273_),
    .ZN(_2274_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5928_ (.A1(_2267_),
    .A2(_2269_),
    .B(_2268_),
    .ZN(_2275_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5929_ (.A1(\r1[5] ),
    .A2(_0377_),
    .ZN(_2276_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5930_ (.A1(\r1[5] ),
    .A2(_0377_),
    .A3(_2275_),
    .ZN(_2277_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5931_ (.A1(net45),
    .A2(_2277_),
    .B(_2274_),
    .C(net34),
    .ZN(_2278_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5932_ (.A1(net13),
    .A2(_2273_),
    .ZN(_2279_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5933_ (.A1(\r1[5] ),
    .A2(net56),
    .ZN(_2280_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5934_ (.A1(\r1[5] ),
    .A2(net56),
    .ZN(_2281_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5935_ (.A1(_2261_),
    .A2(_2262_),
    .B(_2259_),
    .ZN(_2282_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5936_ (.A1(\r1[5] ),
    .A2(net56),
    .A3(_2282_),
    .ZN(_2283_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5937_ (.A1(_2215_),
    .A2(_2283_),
    .B(_2279_),
    .C(net38),
    .ZN(_2284_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5938_ (.A1(_2278_),
    .A2(_2284_),
    .B(net167),
    .ZN(_0093_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5939_ (.A1(_2614_),
    .A2(_2878_),
    .ZN(_2285_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5940_ (.A1(_2614_),
    .A2(_2878_),
    .ZN(_2286_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5941_ (.A1(_2281_),
    .A2(_2282_),
    .B(_2280_),
    .ZN(_2287_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5942_ (.A1(\r1[6] ),
    .A2(_2879_),
    .A3(_2287_),
    .ZN(_2288_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5943_ (.A1(net90),
    .A2(_2614_),
    .B(_2215_),
    .ZN(_2289_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5944_ (.A1(_2214_),
    .A2(_2288_),
    .B(net34),
    .ZN(_2290_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5945_ (.A1(_2614_),
    .A2(_0424_),
    .A3(_0425_),
    .ZN(_2291_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _5946_ (.A1(\r1[5] ),
    .A2(_0377_),
    .B1(_2267_),
    .B2(_2269_),
    .C(_2268_),
    .ZN(_2292_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5947_ (.A1(_2276_),
    .A2(_2292_),
    .Z(_2293_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5948_ (.A1(_2291_),
    .A2(_2293_),
    .ZN(_2294_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5949_ (.A1(_2596_),
    .A2(\r1[6] ),
    .B(net29),
    .ZN(_2295_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5950_ (.A1(net29),
    .A2(_2294_),
    .B(_2295_),
    .ZN(_2296_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5951_ (.A1(_2289_),
    .A2(_2290_),
    .B1(_2296_),
    .B2(net34),
    .ZN(_2297_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5952_ (.A1(net167),
    .A2(_2297_),
    .ZN(_0094_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5953_ (.A1(\r1[7] ),
    .A2(_2876_),
    .ZN(_2298_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5954_ (.A1(\r1[7] ),
    .A2(_2876_),
    .ZN(_2299_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5955_ (.A1(_2286_),
    .A2(_2287_),
    .B(_2285_),
    .ZN(_2300_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5956_ (.A1(\r1[7] ),
    .A2(_2876_),
    .A3(_2300_),
    .ZN(_2301_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5957_ (.A1(net84),
    .A2(\r1[7] ),
    .ZN(_2302_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5958_ (.A1(_2215_),
    .A2(_2302_),
    .ZN(_2303_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5959_ (.A1(_2215_),
    .A2(_2301_),
    .B(_2303_),
    .C(net38),
    .ZN(_2304_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai33_1 _5960_ (.A1(_2614_),
    .A2(_0426_),
    .A3(_0427_),
    .B1(_2276_),
    .B2(_2291_),
    .B3(_2292_),
    .ZN(_2305_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _5961_ (.A1(_2615_),
    .A2(_0476_),
    .A3(_0477_),
    .ZN(_2306_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5962_ (.A1(_0476_),
    .A2(_0477_),
    .B(_2615_),
    .ZN(_2307_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _5963_ (.A1(\r1[7] ),
    .A2(_0478_),
    .A3(_2305_),
    .ZN(_2308_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5964_ (.A1(net45),
    .A2(_2302_),
    .B(net38),
    .ZN(_2309_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5965_ (.A1(net45),
    .A2(_2308_),
    .B(_2309_),
    .ZN(_2310_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5966_ (.A1(_2304_),
    .A2(_2310_),
    .B(net167),
    .ZN(_0095_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5967_ (.A1(\r1[8] ),
    .A2(_0519_),
    .ZN(_2311_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5968_ (.A1(\r1[8] ),
    .A2(_0519_),
    .ZN(_2312_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _5969_ (.A1(net8),
    .A2(_2307_),
    .B(_2306_),
    .ZN(_2313_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5970_ (.A1(_2312_),
    .A2(_2313_),
    .ZN(_2314_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5971_ (.A1(_2312_),
    .A2(_2313_),
    .ZN(_2315_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5972_ (.A1(net29),
    .A2(_2315_),
    .ZN(_2316_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5973_ (.A1(\r1[8] ),
    .A2(_2226_),
    .ZN(_2317_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5974_ (.A1(_2314_),
    .A2(_2316_),
    .B(_2317_),
    .C(net34),
    .ZN(_2318_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5975_ (.A1(_2299_),
    .A2(_2300_),
    .B(_2298_),
    .ZN(_2319_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5976_ (.A1(_2891_),
    .A2(_2319_),
    .ZN(_2320_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5977_ (.A1(_2891_),
    .A2(_2319_),
    .ZN(_2321_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _5978_ (.A1(net84),
    .A2(\r1[8] ),
    .A3(net13),
    .ZN(_2322_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _5979_ (.A1(net13),
    .A2(_2321_),
    .B(_2322_),
    .C(net39),
    .ZN(_2323_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _5980_ (.A1(net169),
    .A2(_2318_),
    .A3(_2323_),
    .Z(_0096_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5981_ (.A1(_2312_),
    .A2(_2313_),
    .B(_2311_),
    .ZN(_2324_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5982_ (.A1(net11),
    .A2(_0518_),
    .B(_0516_),
    .ZN(_2325_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _5983_ (.A1(_2580_),
    .A2(_0319_),
    .B1(_0514_),
    .B2(_2876_),
    .ZN(_2326_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5984_ (.A1(_2581_),
    .A2(_0318_),
    .B(_2582_),
    .ZN(_2327_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _5985_ (.A1(\hvsync_gen.vpos[8] ),
    .A2(_0319_),
    .ZN(_2328_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _5986_ (.A1(_2581_),
    .A2(_2328_),
    .B(_2327_),
    .ZN(_2329_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5987_ (.A1(_2876_),
    .A2(_2329_),
    .ZN(_2330_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5988_ (.A1(_2326_),
    .A2(_2330_),
    .ZN(_2331_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _5989_ (.A1(_2326_),
    .A2(_2330_),
    .Z(_2332_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _5990_ (.I(_2332_),
    .ZN(_2333_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5991_ (.A1(_2325_),
    .A2(_2332_),
    .ZN(_2334_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _5992_ (.A1(\r1[9] ),
    .A2(_2334_),
    .Z(_2335_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5993_ (.A1(\r1[9] ),
    .A2(_2334_),
    .ZN(_2336_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _5994_ (.A1(\r1[9] ),
    .A2(_2334_),
    .Z(_2337_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _5995_ (.A1(_2336_),
    .A2(_2337_),
    .ZN(_2338_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _5996_ (.A1(_2324_),
    .A2(_2338_),
    .ZN(_2339_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _5997_ (.A1(\r1[9] ),
    .A2(_2226_),
    .B1(_2339_),
    .B2(net28),
    .ZN(_2340_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _5998_ (.A1(_2616_),
    .A2(_2876_),
    .B(_2320_),
    .ZN(_2341_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _5999_ (.A1(\r1[9] ),
    .A2(_2214_),
    .A3(_2341_),
    .Z(_2342_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6000_ (.A1(net89),
    .A2(net13),
    .ZN(_2343_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6001_ (.A1(net36),
    .A2(_2343_),
    .ZN(_2344_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6002_ (.A1(_2214_),
    .A2(_2341_),
    .B(\r1[9] ),
    .ZN(_2345_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai32_1 _6003_ (.A1(_2342_),
    .A2(_2344_),
    .A3(_2345_),
    .B1(_2340_),
    .B2(net36),
    .ZN(_2346_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _6004_ (.A1(net169),
    .A2(_2346_),
    .Z(_0097_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6005_ (.A1(_2325_),
    .A2(_2333_),
    .B(_2331_),
    .ZN(_2347_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6006_ (.A1(\hvsync_gen.vpos[7] ),
    .A2(_2328_),
    .ZN(_2348_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6007_ (.A1(_2877_),
    .A2(_2329_),
    .B(_2348_),
    .ZN(_2349_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _6008_ (.A1(_2583_),
    .A2(_2328_),
    .A3(_2349_),
    .ZN(_2350_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6009_ (.A1(_2347_),
    .A2(_2350_),
    .ZN(_2351_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6010_ (.A1(net98),
    .A2(net6),
    .ZN(_2352_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6011_ (.A1(net98),
    .A2(net6),
    .ZN(_2353_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6012_ (.A1(_2324_),
    .A2(_2337_),
    .B(_2335_),
    .ZN(_2354_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _6013_ (.A1(net98),
    .A2(_2342_),
    .Z(_2355_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6014_ (.A1(net98),
    .A2(_2343_),
    .B(_2342_),
    .ZN(_2356_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6015_ (.A1(net82),
    .A2(net98),
    .B(net28),
    .ZN(_2357_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor3_1 _6016_ (.A1(net98),
    .A2(net6),
    .A3(_2354_),
    .Z(_2358_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _6017_ (.A1(net28),
    .A2(_2358_),
    .B(_2357_),
    .C(net35),
    .ZN(_2359_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _6018_ (.A1(net33),
    .A2(_2355_),
    .A3(_2356_),
    .ZN(_2360_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6019_ (.A1(_2359_),
    .A2(_2360_),
    .ZN(_2361_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6020_ (.A1(net164),
    .A2(_2361_),
    .ZN(_0098_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6021_ (.A1(_2353_),
    .A2(_2354_),
    .B(_2352_),
    .ZN(_2362_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6022_ (.A1(\r1[11] ),
    .A2(net6),
    .ZN(_2363_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _6023_ (.I(_2363_),
    .ZN(_2364_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _6024_ (.A1(\r1[11] ),
    .A2(net6),
    .Z(_2365_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6025_ (.A1(_2363_),
    .A2(_2365_),
    .ZN(_2366_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6026_ (.A1(_2362_),
    .A2(_2366_),
    .ZN(_2367_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _6027_ (.A1(\r1[11] ),
    .A2(_2226_),
    .B1(_2367_),
    .B2(net28),
    .ZN(_2368_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6028_ (.A1(net35),
    .A2(_2368_),
    .ZN(_2369_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6029_ (.A1(\r1[11] ),
    .A2(_2343_),
    .B(_2355_),
    .ZN(_2370_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _6030_ (.A1(\r1[11] ),
    .A2(_2355_),
    .Z(_2371_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _6031_ (.A1(net33),
    .A2(_2370_),
    .A3(_2371_),
    .ZN(_2372_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6032_ (.A1(_2369_),
    .A2(_2372_),
    .ZN(_2373_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6033_ (.A1(net164),
    .A2(_2373_),
    .ZN(_0099_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6034_ (.A1(\r1[12] ),
    .A2(net6),
    .ZN(_2374_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6035_ (.A1(\r1[12] ),
    .A2(net6),
    .ZN(_2375_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _6036_ (.A1(_2362_),
    .A2(_2365_),
    .B(_2364_),
    .ZN(_2376_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _6037_ (.A1(_2375_),
    .A2(_2376_),
    .Z(_2377_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6038_ (.A1(_2375_),
    .A2(_2376_),
    .B(net44),
    .ZN(_2378_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _6039_ (.A1(\r1[12] ),
    .A2(_2226_),
    .B1(_2377_),
    .B2(_2378_),
    .C(net35),
    .ZN(_2379_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6040_ (.A1(\r1[12] ),
    .A2(_2343_),
    .B(_2371_),
    .ZN(_2380_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _6041_ (.A1(\r1[12] ),
    .A2(_2371_),
    .Z(_2381_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6042_ (.A1(_2380_),
    .A2(_2381_),
    .B(net35),
    .ZN(_2382_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6043_ (.A1(net169),
    .A2(_2382_),
    .ZN(_2383_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6044_ (.A1(_2379_),
    .A2(_2383_),
    .ZN(_0100_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6045_ (.A1(\r1[13] ),
    .A2(_2226_),
    .ZN(_2384_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6046_ (.A1(\r1[13] ),
    .A2(net6),
    .ZN(_2385_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6047_ (.A1(_2374_),
    .A2(_2377_),
    .B(_2385_),
    .ZN(_2386_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _6048_ (.A1(_2374_),
    .A2(_2377_),
    .A3(_2385_),
    .Z(_2387_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _6049_ (.A1(net44),
    .A2(_2386_),
    .A3(_2387_),
    .B(_2384_),
    .ZN(_2388_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6050_ (.A1(\r1[13] ),
    .A2(_2381_),
    .ZN(_2389_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _6051_ (.I(_2389_),
    .ZN(_2390_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _6052_ (.A1(\r1[13] ),
    .A2(net35),
    .A3(_2343_),
    .ZN(_2391_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6053_ (.A1(net35),
    .A2(_2381_),
    .ZN(_2392_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6054_ (.A1(_2391_),
    .A2(_2392_),
    .ZN(_2393_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _6055_ (.A1(net33),
    .A2(_2388_),
    .B1(_2389_),
    .B2(_2393_),
    .ZN(_2394_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6056_ (.A1(net164),
    .A2(_2394_),
    .ZN(_0101_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6057_ (.A1(\r1[14] ),
    .A2(_2226_),
    .ZN(_2395_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _6058_ (.A1(\r1[14] ),
    .A2(net7),
    .Z(_2396_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6059_ (.A1(\r1[14] ),
    .A2(net7),
    .ZN(_2397_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6060_ (.A1(_2396_),
    .A2(_2397_),
    .ZN(_2398_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6061_ (.A1(\r1[12] ),
    .A2(\r1[13] ),
    .B(net6),
    .ZN(_2399_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _6062_ (.A1(_2375_),
    .A2(_2376_),
    .A3(_2385_),
    .B(_2399_),
    .ZN(_2400_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _6063_ (.A1(_2398_),
    .A2(_2400_),
    .Z(_2401_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6064_ (.A1(_2398_),
    .A2(_2400_),
    .ZN(_2402_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _6065_ (.A1(net44),
    .A2(_2401_),
    .A3(_2402_),
    .B(_2395_),
    .ZN(_2403_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6066_ (.A1(net33),
    .A2(_2403_),
    .ZN(_2404_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6067_ (.A1(\r1[14] ),
    .A2(_2389_),
    .ZN(_2405_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _6068_ (.A1(net36),
    .A2(_2343_),
    .A3(_2405_),
    .ZN(_2406_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6069_ (.A1(_2404_),
    .A2(_2406_),
    .B(net164),
    .ZN(_0102_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _6070_ (.A1(_2396_),
    .A2(_2401_),
    .Z(_2407_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _6071_ (.A1(\r1[15] ),
    .A2(net6),
    .Z(_2408_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6072_ (.A1(_2396_),
    .A2(_2401_),
    .B(_2408_),
    .ZN(_2409_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _6073_ (.A1(_2407_),
    .A2(_2408_),
    .B(_2409_),
    .C(net28),
    .ZN(_2410_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6074_ (.A1(\r1[15] ),
    .A2(_2226_),
    .B(net36),
    .ZN(_2411_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _6075_ (.A1(\r1[14] ),
    .A2(\r1[15] ),
    .A3(_2390_),
    .Z(_2412_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_1 _6076_ (.A1(\r1[15] ),
    .A2(_2343_),
    .B1(_2390_),
    .B2(\r1[14] ),
    .ZN(_2413_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _6077_ (.A1(_2412_),
    .A2(_2413_),
    .Z(_2414_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _6078_ (.A1(_2410_),
    .A2(_2411_),
    .B1(_2414_),
    .B2(net36),
    .C(net164),
    .ZN(_0103_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6079_ (.A1(\r1[16] ),
    .A2(net7),
    .ZN(_2415_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6080_ (.A1(_2618_),
    .A2(net7),
    .ZN(_2416_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6081_ (.A1(_2963_),
    .A2(net7),
    .ZN(_2417_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _6082_ (.I(_2417_),
    .ZN(_2418_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6083_ (.A1(_2398_),
    .A2(_2408_),
    .ZN(_2419_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _6084_ (.A1(_2375_),
    .A2(_2376_),
    .A3(_2385_),
    .A4(_2419_),
    .ZN(_2420_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6085_ (.A1(_2418_),
    .A2(_2420_),
    .ZN(_2421_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6086_ (.A1(_2418_),
    .A2(_2420_),
    .B(_2416_),
    .ZN(_2422_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6087_ (.A1(\r1[16] ),
    .A2(_2412_),
    .ZN(_2423_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6088_ (.A1(net89),
    .A2(net13),
    .B(_2618_),
    .ZN(_2424_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6089_ (.A1(net89),
    .A2(_2618_),
    .B(net44),
    .ZN(_2425_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6090_ (.A1(_2416_),
    .A2(_2421_),
    .ZN(_2426_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _6091_ (.A1(net44),
    .A2(_2426_),
    .B(_2425_),
    .C(net33),
    .ZN(_2427_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _6092_ (.A1(_2412_),
    .A2(_2424_),
    .B(_2423_),
    .C(net35),
    .ZN(_2428_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6093_ (.A1(_2427_),
    .A2(_2428_),
    .B(net164),
    .ZN(_0104_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6094_ (.A1(\r1[17] ),
    .A2(net7),
    .ZN(_2429_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _6095_ (.A1(_2415_),
    .A2(_2422_),
    .A3(_2429_),
    .Z(_2430_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6096_ (.A1(_2415_),
    .A2(_2422_),
    .B(_2429_),
    .ZN(_2431_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or3_1 _6097_ (.A1(net44),
    .A2(_2430_),
    .A3(_2431_),
    .Z(_2432_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6098_ (.A1(\r1[17] ),
    .A2(_2226_),
    .B(net35),
    .ZN(_2433_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _6099_ (.A1(\r1[17] ),
    .A2(_2343_),
    .A3(_2423_),
    .ZN(_2434_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6100_ (.A1(_2069_),
    .A2(_2412_),
    .B(net33),
    .ZN(_2435_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _6101_ (.A1(_2432_),
    .A2(_2433_),
    .B1(_2434_),
    .B2(_2435_),
    .C(net165),
    .ZN(_0105_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _6102_ (.A1(net171),
    .A2(_1912_),
    .ZN(_2436_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 _6103_ (.I(net20),
    .ZN(_2437_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6104_ (.A1(\title_r[0] ),
    .A2(net76),
    .ZN(_2438_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6105_ (.A1(net20),
    .A2(_2438_),
    .ZN(_0106_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6106_ (.A1(\title_r[0] ),
    .A2(_1880_),
    .ZN(_2439_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6107_ (.A1(net62),
    .A2(_2439_),
    .ZN(_2440_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _6108_ (.A1(\title_r[1] ),
    .A2(net62),
    .B1(net47),
    .B2(\hvsync_gen.vpos[0] ),
    .C(_2440_),
    .ZN(_2441_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _6109_ (.A1(_2566_),
    .A2(net46),
    .A3(_2439_),
    .ZN(_2442_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _6110_ (.A1(_2436_),
    .A2(_2441_),
    .A3(_2442_),
    .ZN(_0107_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6111_ (.A1(_1878_),
    .A2(_1883_),
    .B(_1882_),
    .ZN(_2443_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _6112_ (.A1(_1929_),
    .A2(_1930_),
    .A3(_1931_),
    .Z(_2444_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6113_ (.A1(net47),
    .A2(_2443_),
    .ZN(_2445_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _6114_ (.A1(_2752_),
    .A2(_1932_),
    .A3(_2444_),
    .ZN(_2446_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _6115_ (.A1(_1884_),
    .A2(_2445_),
    .B(_2446_),
    .C(net62),
    .ZN(_2447_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _6116_ (.A1(_2542_),
    .A2(net62),
    .B(net20),
    .C(_2447_),
    .ZN(_0108_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _6117_ (.A1(_1877_),
    .A2(_1878_),
    .A3(_1884_),
    .ZN(_2448_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_1 _6118_ (.A1(net46),
    .A2(_1886_),
    .A3(_2448_),
    .ZN(_2449_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _6119_ (.A1(_1932_),
    .A2(_1933_),
    .Z(_2450_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6120_ (.A1(_2751_),
    .A2(_2450_),
    .B(net63),
    .ZN(_2451_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _6121_ (.A1(_2541_),
    .A2(net62),
    .B1(_2449_),
    .B2(_2451_),
    .C(net20),
    .ZN(_0109_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6122_ (.A1(_1934_),
    .A2(_1936_),
    .ZN(_2452_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6123_ (.A1(net46),
    .A2(_1937_),
    .ZN(_2453_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6124_ (.A1(_2452_),
    .A2(_2453_),
    .B(net62),
    .ZN(_2454_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6125_ (.A1(_1887_),
    .A2(_1889_),
    .ZN(_2455_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6126_ (.A1(net46),
    .A2(_2455_),
    .ZN(_2456_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _6127_ (.A1(_2540_),
    .A2(net62),
    .B1(_2454_),
    .B2(_2456_),
    .C(_2436_),
    .ZN(_0110_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6128_ (.A1(_1938_),
    .A2(_1939_),
    .ZN(_2457_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6129_ (.A1(net47),
    .A2(_2457_),
    .ZN(_2458_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6130_ (.A1(_1874_),
    .A2(_1891_),
    .ZN(_2459_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _6131_ (.A1(net47),
    .A2(_2459_),
    .B(_2458_),
    .C(net76),
    .ZN(_2460_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6132_ (.A1(\title_r[5] ),
    .A2(net76),
    .B(_2460_),
    .ZN(_2461_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6133_ (.A1(net20),
    .A2(_2461_),
    .ZN(_0111_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_1 _6134_ (.A1(\title_r[6] ),
    .A2(net156),
    .A3(_1892_),
    .ZN(_2462_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6135_ (.A1(_2752_),
    .A2(_2462_),
    .ZN(_2463_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6136_ (.A1(_1942_),
    .A2(_1944_),
    .ZN(_2464_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6137_ (.A1(_1595_),
    .A2(_1945_),
    .ZN(_2465_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6138_ (.A1(_2464_),
    .A2(_2465_),
    .B(net62),
    .ZN(_2466_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _6139_ (.A1(_2539_),
    .A2(net62),
    .B1(_2463_),
    .B2(_2466_),
    .C(net20),
    .ZN(_0112_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6140_ (.A1(_1946_),
    .A2(_1947_),
    .ZN(_2467_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6141_ (.A1(net47),
    .A2(_2467_),
    .ZN(_2468_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6142_ (.A1(_1869_),
    .A2(_1893_),
    .ZN(_2469_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _6143_ (.A1(net47),
    .A2(_2469_),
    .B(_2468_),
    .C(net76),
    .ZN(_2470_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6144_ (.A1(_2437_),
    .A2(_2470_),
    .ZN(_2471_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6145_ (.A1(_2538_),
    .A2(net63),
    .B(_2471_),
    .ZN(_0113_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6146_ (.A1(_1895_),
    .A2(_1897_),
    .B(net47),
    .ZN(_2472_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6147_ (.A1(_1895_),
    .A2(_1897_),
    .B(_2472_),
    .ZN(_2473_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__mux2_1 _6148_ (.I0(_2538_),
    .I1(_1953_),
    .S(_1957_),
    .Z(_2474_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6149_ (.A1(_1950_),
    .A2(_2474_),
    .ZN(_2475_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _6150_ (.A1(_1950_),
    .A2(_2474_),
    .Z(_2476_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6151_ (.A1(_1594_),
    .A2(_2476_),
    .B(net63),
    .ZN(_2477_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _6152_ (.A1(_2537_),
    .A2(net63),
    .B1(_2473_),
    .B2(_2477_),
    .C(net20),
    .ZN(_0114_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6153_ (.A1(_1953_),
    .A2(_1957_),
    .B(_2475_),
    .ZN(_2478_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or2_1 _6154_ (.A1(_1960_),
    .A2(_2478_),
    .Z(_2479_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6155_ (.A1(_2751_),
    .A2(_2479_),
    .ZN(_2480_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6156_ (.A1(_1960_),
    .A2(_2478_),
    .B(_2480_),
    .ZN(_2481_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6157_ (.A1(_2537_),
    .A2(net152),
    .B(_1898_),
    .ZN(_2482_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6158_ (.A1(_1868_),
    .A2(_2482_),
    .ZN(_2483_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _6159_ (.A1(net46),
    .A2(_2483_),
    .B(_2481_),
    .C(net63),
    .ZN(_2484_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _6160_ (.A1(_2536_),
    .A2(net63),
    .B(net20),
    .C(_2484_),
    .ZN(_0115_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6161_ (.A1(_1899_),
    .A2(_1905_),
    .ZN(_2485_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6162_ (.A1(_1903_),
    .A2(_2485_),
    .ZN(_2486_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6163_ (.A1(_1959_),
    .A2(_2479_),
    .B(_1961_),
    .ZN(_2487_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _6164_ (.A1(_1959_),
    .A2(_1961_),
    .A3(_2479_),
    .Z(_2488_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6165_ (.A1(_2487_),
    .A2(_2488_),
    .B(net47),
    .ZN(_2489_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6166_ (.A1(net63),
    .A2(_2436_),
    .ZN(_2490_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai211_1 _6167_ (.A1(\title_r[10] ),
    .A2(net76),
    .B(_2437_),
    .C(_2489_),
    .ZN(_2491_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6168_ (.A1(_1910_),
    .A2(_2486_),
    .B(_2491_),
    .ZN(_0116_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6169_ (.A1(_1903_),
    .A2(_2485_),
    .B(_1901_),
    .ZN(_2492_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _6170_ (.A1(_1900_),
    .A2(_2492_),
    .Z(_2493_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6171_ (.A1(_1951_),
    .A2(_1955_),
    .B(_2487_),
    .ZN(_2494_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6172_ (.A1(_1964_),
    .A2(_2494_),
    .ZN(_2495_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _6173_ (.A1(\title_r[11] ),
    .A2(net76),
    .B1(net46),
    .B2(_2495_),
    .ZN(_2496_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _6174_ (.A1(_1910_),
    .A2(_2493_),
    .B(_2496_),
    .C(net20),
    .ZN(_0117_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__or3_1 _6175_ (.A1(_1867_),
    .A2(_1904_),
    .A3(_1907_),
    .Z(_2497_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6176_ (.A1(_1908_),
    .A2(_2497_),
    .B(_2751_),
    .ZN(_2498_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6177_ (.A1(\title_r[12] ),
    .A2(_1962_),
    .ZN(_2499_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _6178_ (.A1(\title_r[12] ),
    .A2(net76),
    .B1(net46),
    .B2(_2499_),
    .ZN(_2500_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_1 _6179_ (.A1(net76),
    .A2(_2498_),
    .B(_2500_),
    .C(net20),
    .ZN(_0118_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6180_ (.A1(\title_r[6] ),
    .A2(\title_r[5] ),
    .ZN(_2501_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and4_1 _6181_ (.A1(_2537_),
    .A2(_2538_),
    .A3(_2540_),
    .A4(_2501_),
    .Z(_2502_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_1 _6182_ (.A1(_2534_),
    .A2(_2535_),
    .A3(_2536_),
    .A4(_2502_),
    .ZN(_2503_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6183_ (.A1(\title_r[12] ),
    .A2(_2503_),
    .B(_2565_),
    .ZN(_2504_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _6184_ (.A1(net154),
    .A2(_2750_),
    .A3(_2490_),
    .A4(_2504_),
    .ZN(_2505_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _6185_ (.A1(_1595_),
    .A2(_2436_),
    .ZN(_2506_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6186_ (.A1(_1594_),
    .A2(_2437_),
    .ZN(_2507_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6187_ (.A1(_2505_),
    .A2(_2507_),
    .B(_2592_),
    .ZN(_2508_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6188_ (.A1(_2592_),
    .A2(_2505_),
    .B(_2508_),
    .ZN(_0119_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _6189_ (.A1(\title_r_pixels_in_scanline[1] ),
    .A2(_2508_),
    .Z(_2509_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6190_ (.A1(\title_r_pixels_in_scanline[1] ),
    .A2(_2508_),
    .ZN(_2510_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _6191_ (.A1(_2506_),
    .A2(_2509_),
    .A3(_2510_),
    .ZN(_0120_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6192_ (.A1(\title_r_pixels_in_scanline[2] ),
    .A2(_2509_),
    .ZN(_2511_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6193_ (.A1(_2506_),
    .A2(_2511_),
    .ZN(_0121_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6194_ (.A1(\title_r_pixels_in_scanline[2] ),
    .A2(_2509_),
    .B(\title_r_pixels_in_scanline[3] ),
    .ZN(_2512_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _6195_ (.A1(\title_r_pixels_in_scanline[3] ),
    .A2(\title_r_pixels_in_scanline[2] ),
    .A3(_2509_),
    .Z(_2513_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor3_1 _6196_ (.A1(_2506_),
    .A2(_2512_),
    .A3(_2513_),
    .ZN(_0122_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6197_ (.A1(\title_r_pixels_in_scanline[4] ),
    .A2(_2513_),
    .ZN(_2514_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6198_ (.A1(\title_r_pixels_in_scanline[4] ),
    .A2(_2513_),
    .ZN(_2515_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6199_ (.A1(_2506_),
    .A2(_2515_),
    .ZN(_0123_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xor2_1 _6200_ (.A1(\title_r_pixels_in_scanline[5] ),
    .A2(_2514_),
    .Z(_2516_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6201_ (.A1(_2506_),
    .A2(_2516_),
    .ZN(_0124_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and4_1 _6202_ (.A1(net96),
    .A2(net97),
    .A3(\hvsync_gen.vpos[9] ),
    .A4(_2758_),
    .Z(_2517_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6203_ (.A1(_2757_),
    .A2(_2517_),
    .ZN(_2518_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _6204_ (.A1(net171),
    .A2(_2148_),
    .A3(_2518_),
    .ZN(_2519_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6205_ (.A1(\hvsync_gen.vpos[0] ),
    .A2(_2149_),
    .ZN(_2520_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai21_1 _6206_ (.A1(\hvsync_gen.vpos[0] ),
    .A2(_2519_),
    .B(_2520_),
    .ZN(_0125_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai32_1 _6207_ (.A1(_2758_),
    .A2(_2178_),
    .A3(_2519_),
    .B1(net27),
    .B2(_2577_),
    .ZN(_0126_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6208_ (.A1(net97),
    .A2(_2178_),
    .ZN(_2521_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _6209_ (.A1(_2578_),
    .A2(net27),
    .B1(_2519_),
    .B2(_2521_),
    .ZN(_0127_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6210_ (.A1(net95),
    .A2(_2149_),
    .ZN(_2522_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and3_1 _6211_ (.A1(net95),
    .A2(net97),
    .A3(_2178_),
    .Z(_2523_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _6212_ (.A1(_2179_),
    .A2(_2519_),
    .A3(_2523_),
    .B(_2522_),
    .ZN(_0128_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6213_ (.A1(net94),
    .A2(_2523_),
    .ZN(_2524_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _6214_ (.A1(_2579_),
    .A2(net27),
    .B1(_2519_),
    .B2(_2524_),
    .ZN(_0129_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand2_1 _6215_ (.A1(net93),
    .A2(_2149_),
    .ZN(_2525_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6216_ (.A1(net94),
    .A2(_2523_),
    .B(net93),
    .ZN(_2526_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__and2_1 _6217_ (.A1(_1971_),
    .A2(_2178_),
    .Z(_2527_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai31_1 _6218_ (.A1(_2519_),
    .A2(_2526_),
    .A3(_2527_),
    .B(_2525_),
    .ZN(_0130_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_1 _6219_ (.A1(net91),
    .A2(_2527_),
    .ZN(_2528_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _6220_ (.A1(_2580_),
    .A2(net27),
    .B1(_2519_),
    .B2(_2528_),
    .ZN(_0131_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6221_ (.A1(net92),
    .A2(_2527_),
    .B(\hvsync_gen.vpos[7] ),
    .ZN(_2529_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _6222_ (.A1(_2566_),
    .A2(_2577_),
    .A3(_2581_),
    .A4(_1972_),
    .ZN(_2530_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai32_1 _6223_ (.A1(_2519_),
    .A2(_2529_),
    .A3(_2530_),
    .B1(net27),
    .B2(_2581_),
    .ZN(_0132_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_1 _6224_ (.A1(_2757_),
    .A2(_2517_),
    .B1(_2530_),
    .B2(\hvsync_gen.vpos[8] ),
    .C(net167),
    .ZN(_2531_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nor2_1 _6225_ (.A1(_2149_),
    .A2(_2531_),
    .ZN(_2532_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__nand4_1 _6226_ (.A1(net171),
    .A2(_2148_),
    .A3(_2518_),
    .A4(_2530_),
    .ZN(_2533_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_1 _6227_ (.A1(_2582_),
    .A2(_2533_),
    .B(_2532_),
    .ZN(_0133_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__oai22_1 _6228_ (.A1(_2583_),
    .A2(_2532_),
    .B1(_2533_),
    .B2(_2623_),
    .ZN(_0134_),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 _6229_ (.I(\r2[0] ),
    .Z(\r__t[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6230_ (.D(_0012_),
    .CLK(clknet_leaf_31_clk),
    .Q(\note_freq[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6231_ (.D(_0013_),
    .CLK(clknet_leaf_37_clk),
    .Q(\r2[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6232_ (.D(_0014_),
    .CLK(clknet_leaf_38_clk),
    .Q(\r2[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6233_ (.D(_0015_),
    .CLK(clknet_leaf_37_clk),
    .Q(\r2[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6234_ (.D(_0016_),
    .CLK(clknet_leaf_49_clk),
    .Q(\r2[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6235_ (.D(_0017_),
    .CLK(clknet_leaf_36_clk),
    .Q(\r2[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6236_ (.D(_0018_),
    .CLK(clknet_leaf_35_clk),
    .Q(\r2[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6237_ (.D(_0019_),
    .CLK(clknet_leaf_48_clk),
    .Q(\r2[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6238_ (.D(_0020_),
    .CLK(clknet_leaf_49_clk),
    .Q(\r2[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6239_ (.D(_0021_),
    .CLK(clknet_leaf_49_clk),
    .Q(\r2[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6240_ (.D(_0022_),
    .CLK(clknet_leaf_48_clk),
    .Q(\r2[9] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6241_ (.D(_0023_),
    .CLK(clknet_leaf_48_clk),
    .Q(\r2[10] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6242_ (.D(_0024_),
    .CLK(clknet_leaf_47_clk),
    .Q(\r2[11] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6243_ (.D(_0025_),
    .CLK(clknet_leaf_47_clk),
    .Q(\r2[12] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6244_ (.D(_0026_),
    .CLK(clknet_leaf_46_clk),
    .Q(\r2[13] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6245_ (.D(_0027_),
    .CLK(clknet_leaf_44_clk),
    .Q(\r2[14] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6246_ (.D(_0028_),
    .CLK(clknet_leaf_46_clk),
    .Q(\r2[15] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6247_ (.D(_0029_),
    .CLK(clknet_leaf_45_clk),
    .Q(\r2[16] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6248_ (.D(_0030_),
    .CLK(clknet_leaf_45_clk),
    .Q(\r2[17] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6249_ (.D(_0031_),
    .CLK(clknet_leaf_44_clk),
    .Q(\r2[18] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6250_ (.D(_0032_),
    .CLK(clknet_leaf_39_clk),
    .Q(\note_freq[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6251_ (.D(_0033_),
    .CLK(clknet_leaf_41_clk),
    .Q(\note2_freq[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6252_ (.D(_0034_),
    .CLK(clknet_leaf_1_clk),
    .Q(\title_r[13] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6253_ (.D(_0035_),
    .CLK(clknet_leaf_11_clk),
    .Q(uo_out[0]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6254_ (.D(_0036_),
    .CLK(clknet_leaf_11_clk),
    .Q(uo_out[1]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6255_ (.D(_0037_),
    .CLK(clknet_leaf_11_clk),
    .Q(uo_out[2]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6256_ (.D(_0038_),
    .CLK(clknet_leaf_11_clk),
    .Q(uo_out[4]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6257_ (.D(_0039_),
    .CLK(clknet_leaf_10_clk),
    .Q(uo_out[5]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6258_ (.D(_0040_),
    .CLK(clknet_leaf_11_clk),
    .Q(uo_out[6]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6259_ (.D(_0000_),
    .CLK(clknet_leaf_41_clk),
    .Q(\note2_freq[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6260_ (.D(_0001_),
    .CLK(clknet_leaf_40_clk),
    .Q(\note2_freq[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6261_ (.D(_0002_),
    .CLK(clknet_leaf_38_clk),
    .Q(\note2_freq[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6262_ (.D(_0003_),
    .CLK(clknet_leaf_38_clk),
    .Q(\note2_freq[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6263_ (.D(_0004_),
    .CLK(clknet_leaf_39_clk),
    .Q(\note2_freq[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6264_ (.D(_0041_),
    .CLK(clknet_leaf_41_clk),
    .Q(noise),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6265_ (.D(_0042_),
    .CLK(clknet_leaf_43_clk),
    .Q(\noise_counter[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6266_ (.D(_0043_),
    .CLK(clknet_leaf_41_clk),
    .Q(\noise_counter[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6267_ (.D(_0044_),
    .CLK(clknet_leaf_43_clk),
    .Q(\noise_counter[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6268_ (.D(_0045_),
    .CLK(clknet_leaf_41_clk),
    .Q(\note2_counter[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6269_ (.D(_0046_),
    .CLK(clknet_leaf_40_clk),
    .Q(\note2_counter[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6270_ (.D(_0047_),
    .CLK(clknet_leaf_41_clk),
    .Q(\note2_counter[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6271_ (.D(_0048_),
    .CLK(clknet_leaf_40_clk),
    .Q(\note2_counter[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6272_ (.D(_0049_),
    .CLK(clknet_leaf_40_clk),
    .Q(\note2_counter[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6273_ (.D(_0050_),
    .CLK(clknet_leaf_39_clk),
    .Q(\note2_counter[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6274_ (.D(_0051_),
    .CLK(clknet_leaf_39_clk),
    .Q(\note2_counter[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6275_ (.D(_0052_),
    .CLK(clknet_leaf_39_clk),
    .Q(\note2_counter[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6276_ (.D(_0053_),
    .CLK(clknet_leaf_39_clk),
    .Q(\note2_counter[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6277_ (.D(_0054_),
    .CLK(clknet_leaf_41_clk),
    .Q(note2),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6278_ (.D(_0055_),
    .CLK(clknet_leaf_39_clk),
    .Q(\note_counter[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6279_ (.D(_0056_),
    .CLK(clknet_leaf_39_clk),
    .Q(\note_counter[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6280_ (.D(_0057_),
    .CLK(clknet_leaf_30_clk),
    .Q(\note_counter[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6281_ (.D(_0058_),
    .CLK(clknet_leaf_30_clk),
    .Q(\note_counter[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6282_ (.D(_0059_),
    .CLK(clknet_leaf_30_clk),
    .Q(\note_counter[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6283_ (.D(_0060_),
    .CLK(clknet_leaf_30_clk),
    .Q(\note_counter[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6284_ (.D(_0061_),
    .CLK(clknet_leaf_30_clk),
    .Q(\note_counter[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6285_ (.D(_0062_),
    .CLK(clknet_leaf_30_clk),
    .Q(\note_counter[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6286_ (.D(_0063_),
    .CLK(clknet_leaf_31_clk),
    .Q(note),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6287_ (.D(_0064_),
    .CLK(clknet_leaf_5_clk),
    .Q(\hvsync_gen.hpos[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6288_ (.D(_0065_),
    .CLK(clknet_leaf_6_clk),
    .Q(\hvsync_gen.hpos[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6289_ (.D(_0066_),
    .CLK(clknet_leaf_9_clk),
    .Q(\hvsync_gen.hpos[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6290_ (.D(_0067_),
    .CLK(clknet_leaf_10_clk),
    .Q(\hvsync_gen.hpos[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6291_ (.D(_0068_),
    .CLK(clknet_leaf_10_clk),
    .Q(\hvsync_gen.hpos[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6292_ (.D(_0069_),
    .CLK(clknet_leaf_10_clk),
    .Q(\hvsync_gen.hpos[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6293_ (.D(_0070_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\hvsync_gen.hpos[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6294_ (.D(_0071_),
    .CLK(clknet_leaf_0_clk),
    .Q(\hvsync_gen.hpos[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6295_ (.D(_0072_),
    .CLK(clknet_leaf_0_clk),
    .Q(\hvsync_gen.hpos[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6296_ (.D(_0073_),
    .CLK(clknet_leaf_0_clk),
    .Q(\hvsync_gen.hpos[9] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6297_ (.D(_0074_),
    .CLK(clknet_leaf_10_clk),
    .Q(uo_out[3]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6298_ (.D(_0075_),
    .CLK(clknet_leaf_9_clk),
    .Q(uo_out[7]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6299_ (.D(_0076_),
    .CLK(clknet_leaf_41_clk),
    .Q(\center_y[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6300_ (.D(_0077_),
    .CLK(clknet_leaf_38_clk),
    .Q(\center_x[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6301_ (.D(_0078_),
    .CLK(clknet_leaf_38_clk),
    .Q(\center_x[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6302_ (.D(_0079_),
    .CLK(clknet_leaf_31_clk),
    .Q(\center_x[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6303_ (.D(_0080_),
    .CLK(clknet_leaf_31_clk),
    .Q(\center_x[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6304_ (.D(_0081_),
    .CLK(clknet_leaf_31_clk),
    .Q(\center_x[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6305_ (.D(_0082_),
    .CLK(clknet_leaf_38_clk),
    .Q(\center_x[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6306_ (.D(_0083_),
    .CLK(clknet_leaf_38_clk),
    .Q(\frame_counter[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6307_ (.D(_0084_),
    .CLK(clknet_leaf_15_clk),
    .Q(\frame_counter[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6308_ (.D(_0085_),
    .CLK(clknet_leaf_15_clk),
    .Q(\frame_counter[9] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6309_ (.D(_0086_),
    .CLK(clknet_leaf_50_clk),
    .Q(frame_counter_frac),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6310_ (.D(\r__t[0] ),
    .CLK(clknet_leaf_33_clk),
    .Q(\r[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6311_ (.D(\r__t[1] ),
    .CLK(clknet_leaf_32_clk),
    .Q(\r[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6312_ (.D(\r__t[2] ),
    .CLK(clknet_leaf_32_clk),
    .Q(\r[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6313_ (.D(\r__t[3] ),
    .CLK(clknet_leaf_33_clk),
    .Q(\r[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6314_ (.D(\r__t[4] ),
    .CLK(clknet_leaf_34_clk),
    .Q(\r[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6315_ (.D(\r__t[5] ),
    .CLK(clknet_leaf_34_clk),
    .Q(\r[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6316_ (.D(\r__t[6] ),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\r[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6317_ (.D(\r__t[7] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\r[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6318_ (.D(\r__t[8] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\r[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6319_ (.D(\r__t[9] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\r[9] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6320_ (.D(\r__t[10] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\r[10] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6321_ (.D(\r__t[11] ),
    .CLK(clknet_leaf_15_clk),
    .Q(\r[11] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6322_ (.D(\r__t[12] ),
    .CLK(clknet_leaf_10_clk),
    .Q(\r[12] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6323_ (.D(\r__t[13] ),
    .CLK(clknet_leaf_1_clk),
    .Q(\r[13] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6324_ (.D(\r__t[14] ),
    .CLK(clknet_leaf_1_clk),
    .Q(\r[14] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6325_ (.D(\r__t[15] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\r[15] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6326_ (.D(\r__t[16] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\r[16] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6327_ (.D(\r__t[17] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\r[17] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6328_ (.D(\r__t[18] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\r[18] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6329_ (.D(\r__t[19] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\r[19] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6330_ (.D(net106),
    .CLK(clknet_leaf_26_clk),
    .Q(\pp_x_sq[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6331_ (.D(\pp_x_sq__t[2] ),
    .CLK(clknet_leaf_26_clk),
    .Q(\pp_x_sq[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6332_ (.D(\pp_x_sq__t[3] ),
    .CLK(clknet_leaf_26_clk),
    .Q(\pp_x_sq[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6333_ (.D(\pp_x_sq__t[4] ),
    .CLK(clknet_leaf_26_clk),
    .Q(\pp_x_sq[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6334_ (.D(\pp_x_sq__t[5] ),
    .CLK(clknet_leaf_22_clk),
    .Q(\pp_x_sq[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6335_ (.D(\pp_x_sq__t[6] ),
    .CLK(clknet_leaf_27_clk),
    .Q(\pp_x_sq[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6336_ (.D(\pp_x_sq__t[7] ),
    .CLK(clknet_leaf_27_clk),
    .Q(\pp_x_sq[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6337_ (.D(\pp_x_sq__t[8] ),
    .CLK(clknet_leaf_29_clk),
    .Q(\pp_x_sq[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6338_ (.D(\pp_x_sq__t[9] ),
    .CLK(clknet_leaf_29_clk),
    .Q(\pp_x_sq[9] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6339_ (.D(\pp_x_sq__t[10] ),
    .CLK(clknet_leaf_27_clk),
    .Q(\pp_x_sq[10] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6340_ (.D(\pp_x_sq__t[11] ),
    .CLK(clknet_leaf_27_clk),
    .Q(\pp_x_sq[11] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6341_ (.D(\pp_x_sq__t[12] ),
    .CLK(clknet_leaf_28_clk),
    .Q(\pp_x_sq[12] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6342_ (.D(\pp_x_sq__t[13] ),
    .CLK(clknet_leaf_28_clk),
    .Q(\pp_x_sq[13] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6343_ (.D(\pp_x_sq__t[14] ),
    .CLK(clknet_leaf_28_clk),
    .Q(\pp_x_sq[14] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6344_ (.D(\pp_x_sq__t[15] ),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\pp_x_sq[15] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6345_ (.D(\ppp_y__t[0] ),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\ppp_y[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6346_ (.D(\ppp_y__t[1] ),
    .CLK(clknet_leaf_18_clk),
    .Q(\ppp_y[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6347_ (.D(\ppp_y__t[2] ),
    .CLK(clknet_leaf_17_clk),
    .Q(\ppp_y[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6348_ (.D(\ppp_y__t[3] ),
    .CLK(clknet_leaf_17_clk),
    .Q(\ppp_y[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6349_ (.D(\ppp_y__t[4] ),
    .CLK(clknet_leaf_16_clk),
    .Q(\ppp_y[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6350_ (.D(\ppp_y__t[5] ),
    .CLK(clknet_leaf_16_clk),
    .Q(\ppp_y[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6351_ (.D(\ppp_y__t[6] ),
    .CLK(clknet_leaf_16_clk),
    .Q(\ppp_y[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6352_ (.D(\ppp_y__t[7] ),
    .CLK(clknet_leaf_15_clk),
    .Q(\ppp_y[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6353_ (.D(\dot2[0] ),
    .CLK(clknet_leaf_17_clk),
    .Q(\ppp_x[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6354_ (.D(\dot2[1] ),
    .CLK(clknet_leaf_33_clk),
    .Q(\ppp_x[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6355_ (.D(\dot2[2] ),
    .CLK(clknet_leaf_17_clk),
    .Q(\ppp_x[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6356_ (.D(\dot2[3] ),
    .CLK(clknet_leaf_33_clk),
    .Q(\ppp_x[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6357_ (.D(\dot2[4] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\ppp_x[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6358_ (.D(\dot2[5] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\ppp_x[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6359_ (.D(\dot2[6] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\ppp_x[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6360_ (.D(\dot2[7] ),
    .CLK(clknet_leaf_33_clk),
    .Q(\ppp_x[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6361_ (.D(\p_p__t[0] ),
    .CLK(clknet_leaf_18_clk),
    .Q(\p_p[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6362_ (.D(\p_p__t[1] ),
    .CLK(clknet_leaf_18_clk),
    .Q(\p_p[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6363_ (.D(\p_p__t[2] ),
    .CLK(clknet_leaf_19_clk),
    .Q(\p_p[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6364_ (.D(\p_p__t[3] ),
    .CLK(clknet_leaf_19_clk),
    .Q(\p_p[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6365_ (.D(\p_p__t[4] ),
    .CLK(clknet_leaf_19_clk),
    .Q(\p_p[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6366_ (.D(\p_p__t[5] ),
    .CLK(clknet_leaf_19_clk),
    .Q(\p_p[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6367_ (.D(\p_p__t[6] ),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\p_p[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6368_ (.D(\p_p__t[7] ),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\p_p[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6369_ (.D(\dot__t[0] ),
    .CLK(clknet_leaf_22_clk),
    .Q(\dot[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6370_ (.D(\dot__t[1] ),
    .CLK(clknet_leaf_22_clk),
    .Q(\dot[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6371_ (.D(\dot__t[2] ),
    .CLK(clknet_leaf_22_clk),
    .Q(\dot[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6372_ (.D(\dot__t[3] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\dot[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6373_ (.D(\dot__t[4] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\dot[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6374_ (.D(\dot__t[5] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\dot[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6375_ (.D(\dot__t[6] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\dot[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6376_ (.D(\dot__t[7] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\dot[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 _6377_ (.D(_0087_),
    .CLK(clknet_leaf_11_clk),
    .Q(uio_out[7]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6378_ (.D(_0088_),
    .CLK(clknet_leaf_38_clk),
    .Q(\r1[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6379_ (.D(_0089_),
    .CLK(clknet_leaf_38_clk),
    .Q(\r1[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6380_ (.D(_0090_),
    .CLK(clknet_leaf_36_clk),
    .Q(\r1[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6381_ (.D(_0091_),
    .CLK(clknet_leaf_35_clk),
    .Q(\r1[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6382_ (.D(_0092_),
    .CLK(clknet_leaf_35_clk),
    .Q(\r1[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6383_ (.D(_0093_),
    .CLK(clknet_leaf_50_clk),
    .Q(\r1[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6384_ (.D(_0094_),
    .CLK(clknet_leaf_15_clk),
    .Q(\r1[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6385_ (.D(_0095_),
    .CLK(clknet_leaf_50_clk),
    .Q(\r1[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6386_ (.D(_0096_),
    .CLK(clknet_leaf_37_clk),
    .Q(\r1[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6387_ (.D(_0097_),
    .CLK(clknet_leaf_42_clk),
    .Q(\r1[9] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6388_ (.D(_0098_),
    .CLK(clknet_leaf_42_clk),
    .Q(\r1[10] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6389_ (.D(_0099_),
    .CLK(clknet_leaf_44_clk),
    .Q(\r1[11] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6390_ (.D(_0100_),
    .CLK(clknet_leaf_44_clk),
    .Q(\r1[12] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6391_ (.D(_0101_),
    .CLK(clknet_leaf_43_clk),
    .Q(\r1[13] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6392_ (.D(_0102_),
    .CLK(clknet_leaf_43_clk),
    .Q(\r1[14] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6393_ (.D(_0103_),
    .CLK(clknet_leaf_43_clk),
    .Q(\r1[15] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6394_ (.D(_0104_),
    .CLK(clknet_leaf_41_clk),
    .Q(\r1[16] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6395_ (.D(_0105_),
    .CLK(clknet_leaf_41_clk),
    .Q(\r1[17] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6396_ (.D(_0106_),
    .CLK(clknet_leaf_6_clk),
    .Q(\title_r[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6397_ (.D(_0107_),
    .CLK(clknet_leaf_5_clk),
    .Q(\title_r[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6398_ (.D(_0108_),
    .CLK(clknet_leaf_8_clk),
    .Q(\title_r[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6399_ (.D(_0109_),
    .CLK(clknet_leaf_8_clk),
    .Q(\title_r[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6400_ (.D(_0110_),
    .CLK(clknet_leaf_7_clk),
    .Q(\title_r[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6401_ (.D(_0111_),
    .CLK(clknet_leaf_7_clk),
    .Q(\title_r[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6402_ (.D(_0112_),
    .CLK(clknet_leaf_7_clk),
    .Q(\title_r[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6403_ (.D(_0113_),
    .CLK(clknet_leaf_4_clk),
    .Q(\title_r[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6404_ (.D(_0114_),
    .CLK(clknet_leaf_3_clk),
    .Q(\title_r[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6405_ (.D(_0115_),
    .CLK(clknet_leaf_2_clk),
    .Q(\title_r[9] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6406_ (.D(_0116_),
    .CLK(clknet_leaf_2_clk),
    .Q(\title_r[10] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6407_ (.D(_0117_),
    .CLK(clknet_leaf_47_clk),
    .Q(\title_r[11] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6408_ (.D(_0118_),
    .CLK(clknet_leaf_1_clk),
    .Q(\title_r[12] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6409_ (.D(_0119_),
    .CLK(clknet_leaf_4_clk),
    .Q(\title_r_pixels_in_scanline[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6410_ (.D(_0120_),
    .CLK(clknet_leaf_9_clk),
    .Q(\title_r_pixels_in_scanline[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6411_ (.D(_0121_),
    .CLK(clknet_leaf_8_clk),
    .Q(\title_r_pixels_in_scanline[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6412_ (.D(_0122_),
    .CLK(clknet_leaf_9_clk),
    .Q(\title_r_pixels_in_scanline[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6413_ (.D(_0123_),
    .CLK(clknet_leaf_9_clk),
    .Q(\title_r_pixels_in_scanline[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6414_ (.D(_0124_),
    .CLK(clknet_leaf_9_clk),
    .Q(\title_r_pixels_in_scanline[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6415_ (.D(_0010_),
    .CLK(clknet_leaf_9_clk),
    .Q(hsync),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6416_ (.D(_0125_),
    .CLK(clknet_leaf_5_clk),
    .Q(\hvsync_gen.vpos[0] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 _6417_ (.D(_0126_),
    .CLK(clknet_leaf_5_clk),
    .Q(\hvsync_gen.vpos[1] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6418_ (.D(_0127_),
    .CLK(clknet_leaf_5_clk),
    .Q(\hvsync_gen.vpos[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6419_ (.D(_0128_),
    .CLK(clknet_leaf_4_clk),
    .Q(\hvsync_gen.vpos[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6420_ (.D(_0129_),
    .CLK(clknet_leaf_1_clk),
    .Q(\hvsync_gen.vpos[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6421_ (.D(_0130_),
    .CLK(clknet_leaf_3_clk),
    .Q(\hvsync_gen.vpos[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6422_ (.D(_0131_),
    .CLK(clknet_leaf_3_clk),
    .Q(\hvsync_gen.vpos[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6423_ (.D(_0132_),
    .CLK(clknet_leaf_5_clk),
    .Q(\hvsync_gen.vpos[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6424_ (.D(_0133_),
    .CLK(clknet_leaf_1_clk),
    .Q(\hvsync_gen.vpos[8] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6425_ (.D(_0134_),
    .CLK(clknet_leaf_1_clk),
    .Q(\hvsync_gen.vpos[9] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6426_ (.D(_0011_),
    .CLK(clknet_leaf_1_clk),
    .Q(\hvsync_gen.vsync ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6427_ (.D(_0005_),
    .CLK(clknet_leaf_31_clk),
    .Q(\note_freq[2] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6428_ (.D(_0006_),
    .CLK(clknet_leaf_31_clk),
    .Q(\note_freq[4] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6429_ (.D(_0007_),
    .CLK(clknet_leaf_31_clk),
    .Q(\note_freq[5] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6430_ (.D(_0008_),
    .CLK(clknet_leaf_31_clk),
    .Q(\note_freq[6] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6431_ (.D(_0009_),
    .CLK(clknet_leaf_31_clk),
    .Q(\note_freq[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6432_ (.D(_0135_),
    .CLK(clknet_leaf_38_clk),
    .Q(\note2_freq[7] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dffq_1 _6433_ (.D(_0136_),
    .CLK(clknet_leaf_39_clk),
    .Q(\note2_freq[3] ),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__tieh tt_um_rejunity_vga_test01_174 (.Z(net174),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__tieh tt_um_rejunity_vga_test01_175 (.Z(net175),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__tieh tt_um_rejunity_vga_test01_176 (.Z(net176),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__tieh tt_um_rejunity_vga_test01_177 (.Z(net177),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__tieh tt_um_rejunity_vga_test01_178 (.Z(net178),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__tieh tt_um_rejunity_vga_test01_179 (.Z(net179),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__tieh tt_um_rejunity_vga_test01_180 (.Z(net180),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_0_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 _6442_ (.I(uio_out[7]),
    .Z(uio_out[0]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 _6443_ (.I(uio_out[7]),
    .Z(uio_out[1]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 _6444_ (.I(uio_out[7]),
    .Z(uio_out[2]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 _6445_ (.I(uio_out[7]),
    .Z(uio_out[3]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 _6446_ (.I(uio_out[7]),
    .Z(uio_out[4]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 _6447_ (.I(uio_out[7]),
    .Z(uio_out[5]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 _6448_ (.I(uio_out[7]),
    .Z(uio_out[6]),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_62 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_63 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_64 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_65 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_66 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_67 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_68 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_69 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_70 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_71 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_72 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_73 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_74 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_75 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_76 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_77 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_78 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_79 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_80 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_81 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_82 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_83 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_84 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_85 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_86 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_87 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_88 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_89 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_90 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_91 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_92 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_93 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_94 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_95 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_96 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_97 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_98 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_99 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_100 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_101 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_102 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_103 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_104 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_105 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_106 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_107 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_108 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_109 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_110 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_111 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_112 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_113 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_114 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_115 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_116 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_117 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_118 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_119 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_120 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_121 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_122 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_123 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_124 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_125 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_126 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_127 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_128 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_129 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_130 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_131 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_132 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_133 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_134 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_135 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_136 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_137 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_138 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_139 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_140 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_141 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_142 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_143 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_144 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_145 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_146 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_147 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_148 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_149 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_150 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_151 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_152 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_153 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_154 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_155 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_156 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_157 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_158 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_159 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_160 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_161 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_162 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_163 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_164 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_165 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_166 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_167 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_168 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_169 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_170 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_171 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_172 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_173 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_174 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_175 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_176 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_177 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_178 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_179 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_180 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_181 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_182 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_183 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_184 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_185 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_186 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_187 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_188 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_189 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_190 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_191 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_192 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_193 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_194 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_195 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_196 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_197 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_198 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_199 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_200 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_201 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_202 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_203 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_204 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_205 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_206 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_207 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_208 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_209 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_210 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_211 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_212 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_213 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_214 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_215 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_216 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_217 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_218 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_219 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_220 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_221 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_222 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_223 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_224 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_225 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_226 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_227 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_228 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_229 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_230 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_231 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_232 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_233 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_234 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_235 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_236 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_237 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_238 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_239 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_240 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_241 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_242 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_243 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_244 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_245 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_246 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_247 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_248 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_249 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_250 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_251 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_252 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_253 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_254 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_255 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_256 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_257 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_258 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_259 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_260 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_261 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_262 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_263 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_264 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_265 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_266 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_267 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_268 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_269 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_270 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_271 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_272 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_273 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_274 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_275 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_276 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_277 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_278 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_279 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_280 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_281 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_282 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_283 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_284 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_285 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_286 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_287 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_288 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_289 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_290 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_291 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_292 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_293 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_294 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_295 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_296 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_297 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_298 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_299 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_300 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_301 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_302 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_303 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_304 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_305 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_306 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_307 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_308 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_309 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_310 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_311 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_312 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_313 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_314 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_315 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_316 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_317 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_318 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_319 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_320 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_321 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_322 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_323 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_324 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_325 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_326 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_327 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_328 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_329 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_330 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_331 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_332 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_333 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_334 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_335 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_336 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_337 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_338 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_339 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_340 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_341 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_342 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_343 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_344 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_345 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_346 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_347 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_348 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_349 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_350 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_351 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_352 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_353 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_354 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_355 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_356 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_357 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_358 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_359 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_360 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_361 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_362 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_363 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_364 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_365 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_366 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_367 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_368 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_369 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_370 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_371 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_372 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_373 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_374 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_375 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_376 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_377 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_378 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_379 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_380 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_381 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_382 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_383 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_384 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_385 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_386 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_387 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_388 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_389 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_390 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_391 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_392 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_393 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_394 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_395 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_396 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_397 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_398 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_399 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_400 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_401 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_402 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_403 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_404 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_405 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_406 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_407 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_408 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_409 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_410 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_411 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_412 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_413 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_414 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_415 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_416 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_417 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_418 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_419 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_420 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_421 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_422 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_423 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_424 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_425 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_426 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_427 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_428 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_429 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_430 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_431 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_432 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_433 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_434 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_435 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_436 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_437 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_438 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_439 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_440 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_441 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_442 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_443 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_444 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_445 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_446 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_447 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_448 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_449 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_450 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_451 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_452 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_453 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_454 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_455 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_456 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_457 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_458 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_459 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_460 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_461 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_462 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_463 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_464 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_465 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_466 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_467 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_468 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_469 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_470 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_471 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_472 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_473 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_474 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_475 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_476 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_477 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_478 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_479 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_480 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_481 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_482 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_483 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_484 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_485 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_486 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_487 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_488 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_489 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_490 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_491 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_492 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_493 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_494 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_495 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_496 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_497 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_498 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_499 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_500 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_501 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_502 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_503 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_504 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_505 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_506 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_507 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_508 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_509 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_510 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_511 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_512 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_513 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_514 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_515 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_516 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_517 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_518 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_519 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_520 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_521 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_522 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_523 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_524 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_525 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_526 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_527 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_528 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_529 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_530 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_531 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_532 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_533 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_534 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_535 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_536 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_537 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_538 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_539 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_540 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_541 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_542 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_543 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_544 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_545 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_546 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_547 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_548 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_549 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_550 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_551 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_552 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_553 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_554 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_555 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_556 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_557 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_558 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_559 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_560 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_561 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_562 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_563 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_564 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_565 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_566 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_567 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_568 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_569 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_570 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_571 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_572 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_573 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_574 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_575 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_576 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_577 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_578 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_579 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_580 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_581 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_582 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_583 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_584 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_585 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_586 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_587 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_588 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_589 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_590 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_591 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_592 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_593 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_594 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_595 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_596 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_597 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_598 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_599 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_600 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_601 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_602 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_603 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_604 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_605 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_606 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_607 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_608 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_609 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_610 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_611 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_612 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_613 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_614 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_615 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_616 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_617 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_618 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_619 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_620 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_621 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_622 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_623 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_624 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_625 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_626 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_627 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_628 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_629 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_630 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_631 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_632 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_633 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_634 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_635 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_636 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_637 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_638 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_639 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_640 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_641 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_642 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_643 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_644 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_645 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_646 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_647 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_648 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_649 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_650 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_651 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_652 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_653 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_654 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_655 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_656 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_657 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_658 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_659 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_660 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_661 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_662 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_663 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_664 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_665 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_666 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_667 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_668 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_669 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_670 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_671 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_672 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_673 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_674 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_675 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_676 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_677 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_678 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_679 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_680 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_681 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_682 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_683 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_684 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_685 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_686 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_687 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_688 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_689 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_690 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_691 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_692 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_693 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_694 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_695 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_696 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_697 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_698 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_699 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_700 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_701 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_702 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_703 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_704 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_705 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_706 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_707 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_708 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_709 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_710 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_711 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_712 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_713 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_714 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_715 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_716 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_717 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_718 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_719 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_720 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_721 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_722 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_723 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_724 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_725 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_726 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_727 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_728 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_729 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_730 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_731 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_732 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_733 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_734 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_735 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_736 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_737 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_738 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_739 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_740 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_741 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_742 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_743 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_744 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_745 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_746 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_747 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_748 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_749 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_750 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_751 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_752 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_753 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_754 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_755 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_756 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_757 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_758 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_759 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_760 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_761 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_762 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_763 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_764 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_765 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_766 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_767 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_768 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_769 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_770 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_771 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_772 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_773 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_774 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_775 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_776 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_777 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_778 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_779 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_780 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_781 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_782 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_783 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_784 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_785 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_786 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_787 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_788 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_789 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_790 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_791 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_792 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_793 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_794 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_795 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_796 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_797 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_798 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_799 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_800 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_801 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_802 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_803 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_804 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_805 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_806 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_807 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_808 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_809 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_810 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_811 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_812 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_813 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_814 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_815 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_816 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_817 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_818 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_819 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_820 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_821 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_822 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_823 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_824 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_825 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_826 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_827 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_828 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_829 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_830 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_831 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_832 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_833 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_834 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_835 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_836 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_837 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_838 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_839 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_840 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_841 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_842 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_843 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_844 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_845 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_846 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_847 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_848 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_849 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_850 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_851 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_852 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_853 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_854 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_855 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_856 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_857 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_858 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_859 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_860 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_861 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_862 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_863 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_864 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_865 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_866 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_867 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_868 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_869 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_870 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_871 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_872 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_873 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_874 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_875 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_876 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_877 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_878 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_879 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_880 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_881 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_882 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_883 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_884 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_885 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_886 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_887 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_888 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_889 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_890 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_891 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_892 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_893 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_894 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_895 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_896 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_897 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_898 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_899 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_900 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_901 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_902 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_903 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_904 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_905 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_906 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_907 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_908 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_909 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_910 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_911 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_912 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_913 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_914 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_915 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_916 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_917 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_918 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_919 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_920 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_921 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_922 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_923 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_924 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_925 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_926 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_927 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_928 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_929 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_930 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_931 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_932 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_933 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_934 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_935 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_936 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_937 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_938 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_939 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_940 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_941 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_942 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_943 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_944 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_945 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_946 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_947 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_948 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_949 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_950 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_951 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_952 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_953 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_954 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_955 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_956 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_957 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_958 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_959 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_960 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_961 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_962 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_963 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_964 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_965 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_966 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_967 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_968 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_969 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_970 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_971 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_972 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_973 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_974 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_975 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_976 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_977 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_978 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_979 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_980 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_981 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_982 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_983 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_984 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_985 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_986 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_987 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_988 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_989 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_990 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_991 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_992 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_993 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_994 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_995 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_996 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_997 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_998 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_999 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1000 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1001 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1002 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1003 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1004 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1005 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1006 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1007 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1008 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1009 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1010 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1011 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1012 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1013 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1014 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1015 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_1016 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1017 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1018 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1019 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1020 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1021 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1022 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1023 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1024 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1025 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1026 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1027 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1028 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1029 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1030 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1031 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1032 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1033 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_1034 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1035 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1036 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1037 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1038 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1039 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1040 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1041 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1042 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1043 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1044 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1045 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1046 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1047 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1048 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1049 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1050 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_1051 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1052 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1053 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1054 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1055 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1056 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1057 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1058 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1059 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1060 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1061 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1062 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1063 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1064 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1065 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1066 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1067 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1068 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_1069 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1070 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1071 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1072 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1073 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1074 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1075 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1076 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1077 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1078 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1079 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1080 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1081 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1082 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1083 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1084 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1085 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_1086 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1087 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1088 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1089 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1090 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1091 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1092 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1093 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1094 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1095 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1096 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1097 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1098 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1099 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1100 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1101 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1102 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1103 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_1104 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1105 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1106 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1107 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1108 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1109 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1110 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1111 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1112 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1113 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1114 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1115 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1116 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1117 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1118 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1119 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1120 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_1121 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1122 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1123 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1124 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1125 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1126 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1127 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1128 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1129 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1130 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1131 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1132 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1133 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1134 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1135 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1136 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1137 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1138 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_1139 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1140 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1141 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1142 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1143 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1144 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1145 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1146 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1147 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1148 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1149 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1150 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1151 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1152 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1153 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1154 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1155 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_1156 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1157 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1158 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1159 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1160 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1161 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1162 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1163 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1164 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1165 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1166 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1167 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1168 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1169 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1170 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1171 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1172 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1173 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_1174 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1175 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1176 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1177 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1178 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1179 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1180 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1181 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1182 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1183 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1184 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1185 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1186 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1187 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1188 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1189 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1190 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_1191 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1192 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1193 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1194 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1195 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1196 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1197 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1198 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1199 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1200 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1201 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1202 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1203 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1204 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1205 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1206 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1207 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1208 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_1209 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1210 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1211 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1212 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1213 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1214 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1215 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1216 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1217 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1218 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1219 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1220 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1221 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1222 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1223 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1224 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1225 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1226 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1227 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1228 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1229 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1230 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1231 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1232 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1233 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1234 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1235 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1236 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1237 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1238 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1239 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1240 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1241 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1242 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1243 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1244 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_1245 (.VDD(VPWR),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_1 input1 (.I(rst_n),
    .Z(net1),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_1 max_cap2 (.I(_2976_),
    .Z(net2),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_1 wire3 (.I(_0466_),
    .Z(net3),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_1 max_cap4 (.I(_0914_),
    .Z(net4),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_1 max_cap5 (.I(_2940_),
    .Z(net5),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout6 (.I(_2351_),
    .Z(net6),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout7 (.I(_2351_),
    .Z(net7),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_1 max_cap8 (.I(_2305_),
    .Z(net8),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_1 max_cap9 (.I(net10),
    .Z(net9),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_1 wire10 (.I(_0888_),
    .Z(net10),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_1 wire11 (.I(_0510_),
    .Z(net11),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 wire12 (.I(_0428_),
    .Z(net12),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout13 (.I(_2215_),
    .Z(net13),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout14 (.I(net15),
    .Z(net14),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout15 (.I(_1744_),
    .Z(net15),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_1 max_cap16 (.I(_0873_),
    .Z(net16),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 max_cap17 (.I(_0328_),
    .Z(net17),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 max_cap18 (.I(_0282_),
    .Z(net18),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 max_cap19 (.I(_0223_),
    .Z(net19),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout20 (.I(_2436_),
    .Z(net20),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout21 (.I(_1603_),
    .Z(net21),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout22 (.I(_1589_),
    .Z(net22),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout23 (.I(net25),
    .Z(net23),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout24 (.I(net25),
    .Z(net24),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 wire25 (.I(_1588_),
    .Z(net25),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 max_cap26 (.I(_0231_),
    .Z(net26),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout27 (.I(_2150_),
    .Z(net27),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout28 (.I(_1759_),
    .Z(net28),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout29 (.I(_1759_),
    .Z(net29),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout30 (.I(net31),
    .Z(net30),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout31 (.I(_1610_),
    .Z(net31),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout32 (.I(_1609_),
    .Z(net32),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout33 (.I(_1602_),
    .Z(net33),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout34 (.I(_1602_),
    .Z(net34),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout35 (.I(net37),
    .Z(net35),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 fanout36 (.I(net37),
    .Z(net36),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout37 (.I(_1601_),
    .Z(net37),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout38 (.I(net39),
    .Z(net38),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout39 (.I(_1601_),
    .Z(net39),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout40 (.I(_1597_),
    .Z(net40),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 fanout41 (.I(_1597_),
    .Z(net41),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout42 (.I(_1596_),
    .Z(net42),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 max_cap43 (.I(_2687_),
    .Z(net43),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout44 (.I(net45),
    .Z(net44),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout45 (.I(_1760_),
    .Z(net45),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout46 (.I(_1595_),
    .Z(net46),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout47 (.I(_1594_),
    .Z(net47),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout48 (.I(_0591_),
    .Z(net48),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout49 (.I(_0591_),
    .Z(net49),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout50 (.I(_0590_),
    .Z(net50),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout51 (.I(net53),
    .Z(net51),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout52 (.I(_0559_),
    .Z(net52),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 fanout53 (.I(_0559_),
    .Z(net53),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout54 (.I(_0248_),
    .Z(net54),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout55 (.I(_0226_),
    .Z(net55),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout56 (.I(_2862_),
    .Z(net56),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout57 (.I(_2861_),
    .Z(net57),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout58 (.I(_2754_),
    .Z(net58),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout59 (.I(_2753_),
    .Z(net59),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout60 (.I(_2639_),
    .Z(net60),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 fanout61 (.I(_2639_),
    .Z(net61),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout62 (.I(net63),
    .Z(net62),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout63 (.I(_2627_),
    .Z(net63),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout64 (.I(_0563_),
    .Z(net64),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout65 (.I(_0563_),
    .Z(net65),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout66 (.I(_0561_),
    .Z(net66),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout67 (.I(_0561_),
    .Z(net67),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout68 (.I(_0543_),
    .Z(net68),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout69 (.I(_0543_),
    .Z(net69),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout70 (.I(net71),
    .Z(net70),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout71 (.I(_0234_),
    .Z(net71),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_1 max_cap72 (.I(_3009_),
    .Z(net72),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 max_cap73 (.I(_2989_),
    .Z(net73),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout74 (.I(net75),
    .Z(net74),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout75 (.I(_2778_),
    .Z(net75),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 wire76 (.I(_2626_),
    .Z(net76),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout77 (.I(net78),
    .Z(net77),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout78 (.I(_0539_),
    .Z(net78),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 fanout79 (.I(_0539_),
    .Z(net79),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 fanout80 (.I(_0233_),
    .Z(net80),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 max_cap81 (.I(_2631_),
    .Z(net81),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout82 (.I(_2596_),
    .Z(net82),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 fanout83 (.I(_2596_),
    .Z(net83),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout84 (.I(_2596_),
    .Z(net84),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout85 (.I(net86),
    .Z(net85),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout86 (.I(_2547_),
    .Z(net86),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 fanout87 (.I(_2547_),
    .Z(net87),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 fanout88 (.I(_2546_),
    .Z(net88),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 fanout89 (.I(\hvsync_gen.vsync ),
    .Z(net89),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout90 (.I(\hvsync_gen.vsync ),
    .Z(net90),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout91 (.I(net92),
    .Z(net91),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout92 (.I(\hvsync_gen.vpos[6] ),
    .Z(net92),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout93 (.I(\hvsync_gen.vpos[5] ),
    .Z(net93),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout94 (.I(\hvsync_gen.vpos[4] ),
    .Z(net94),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout95 (.I(net96),
    .Z(net95),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout96 (.I(\hvsync_gen.vpos[3] ),
    .Z(net96),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout97 (.I(\hvsync_gen.vpos[2] ),
    .Z(net97),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout98 (.I(\r1[10] ),
    .Z(net98),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout99 (.I(\dot[7] ),
    .Z(net99),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout100 (.I(net102),
    .Z(net100),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 fanout101 (.I(net102),
    .Z(net101),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout102 (.I(\dot[6] ),
    .Z(net102),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout103 (.I(\dot[5] ),
    .Z(net103),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout104 (.I(\dot[2] ),
    .Z(net104),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout105 (.I(\dot[1] ),
    .Z(net105),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout106 (.I(\dot[0] ),
    .Z(net106),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout107 (.I(\r[12] ),
    .Z(net107),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout108 (.I(\r[3] ),
    .Z(net108),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout109 (.I(\r[2] ),
    .Z(net109),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout110 (.I(\r[1] ),
    .Z(net110),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 fanout111 (.I(\frame_counter[9] ),
    .Z(net111),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 fanout112 (.I(\center_x[5] ),
    .Z(net112),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 fanout113 (.I(\center_x[5] ),
    .Z(net113),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout114 (.I(net115),
    .Z(net114),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout115 (.I(\center_x[5] ),
    .Z(net115),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout116 (.I(net117),
    .Z(net116),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout117 (.I(net118),
    .Z(net117),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout118 (.I(net121),
    .Z(net118),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout119 (.I(net120),
    .Z(net119),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout120 (.I(net121),
    .Z(net120),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout121 (.I(\center_x[4] ),
    .Z(net121),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout122 (.I(net123),
    .Z(net122),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout123 (.I(\center_x[3] ),
    .Z(net123),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout124 (.I(net125),
    .Z(net124),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 fanout125 (.I(\center_x[3] ),
    .Z(net125),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout126 (.I(net127),
    .Z(net126),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout127 (.I(\center_x[2] ),
    .Z(net127),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout128 (.I(net129),
    .Z(net128),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout129 (.I(\center_x[2] ),
    .Z(net129),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout130 (.I(net135),
    .Z(net130),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout131 (.I(net135),
    .Z(net131),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout132 (.I(net134),
    .Z(net132),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout133 (.I(net134),
    .Z(net133),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout134 (.I(net135),
    .Z(net134),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout135 (.I(\center_x[1] ),
    .Z(net135),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout136 (.I(net137),
    .Z(net136),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout137 (.I(net142),
    .Z(net137),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout138 (.I(net140),
    .Z(net138),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout139 (.I(net140),
    .Z(net139),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 fanout140 (.I(net141),
    .Z(net140),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout141 (.I(net142),
    .Z(net141),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout142 (.I(\center_x[0] ),
    .Z(net142),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout143 (.I(net144),
    .Z(net143),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout144 (.I(net151),
    .Z(net144),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout145 (.I(net146),
    .Z(net145),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout146 (.I(net147),
    .Z(net146),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout147 (.I(net150),
    .Z(net147),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout148 (.I(net149),
    .Z(net148),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 fanout149 (.I(net150),
    .Z(net149),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout150 (.I(net151),
    .Z(net150),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout151 (.I(\center_y[0] ),
    .Z(net151),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout152 (.I(net154),
    .Z(net152),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout153 (.I(net154),
    .Z(net153),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout154 (.I(\hvsync_gen.hpos[6] ),
    .Z(net154),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout155 (.I(net156),
    .Z(net155),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout156 (.I(\hvsync_gen.hpos[5] ),
    .Z(net156),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout157 (.I(net159),
    .Z(net157),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 fanout158 (.I(net159),
    .Z(net158),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout159 (.I(\hvsync_gen.hpos[4] ),
    .Z(net159),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout160 (.I(net161),
    .Z(net160),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 fanout161 (.I(\hvsync_gen.hpos[3] ),
    .Z(net161),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 fanout162 (.I(\hvsync_gen.hpos[2] ),
    .Z(net162),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_1 fanout163 (.I(\hvsync_gen.hpos[2] ),
    .Z(net163),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout164 (.I(net165),
    .Z(net164),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout165 (.I(net168),
    .Z(net165),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout166 (.I(net168),
    .Z(net166),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout167 (.I(net168),
    .Z(net167),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 fanout168 (.I(_2584_),
    .Z(net168),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout169 (.I(net170),
    .Z(net169),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 fanout170 (.I(net172),
    .Z(net170),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 fanout171 (.I(net172),
    .Z(net171),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 fanout172 (.I(net1),
    .Z(net172),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__tieh tt_um_rejunity_vga_test01_173 (.Z(net173),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_1_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_1_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_2_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_3_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_3_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_4_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_4_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_5_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_5_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_6_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_6_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_7_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_8_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_8_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_9_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_9_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_10_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_10_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_11_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_11_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_15_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_15_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_16_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_16_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_17_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_17_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_18_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_18_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_19_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_19_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_21_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_21_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_22_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_22_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_23_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_23_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_26_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_26_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_27_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_27_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_28_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_28_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_29_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_29_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_30_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_30_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_31_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_32_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_32_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_33_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_33_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_34_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_34_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_35_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_35_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_36_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_36_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_37_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_37_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_38_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_38_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_39_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_39_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_40_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_40_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_41_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_41_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_42_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_42_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_43_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_43_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_44_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_44_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_45_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_45_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_46_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_46_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_47_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_47_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_48_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_48_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_49_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_49_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clkbuf_leaf_50_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_50_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload0 (.I(clknet_2_1__leaf_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload1 (.I(clknet_2_2__leaf_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload2 (.I(clknet_2_3__leaf_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload3 (.I(clknet_leaf_35_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload4 (.I(clknet_leaf_36_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload5 (.I(clknet_leaf_37_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload6 (.I(clknet_leaf_39_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload7 (.I(clknet_leaf_40_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload8 (.I(clknet_leaf_41_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload9 (.I(clknet_leaf_42_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload10 (.I(clknet_leaf_43_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload11 (.I(clknet_leaf_44_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload12 (.I(clknet_leaf_45_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload13 (.I(clknet_leaf_46_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload14 (.I(clknet_leaf_48_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload15 (.I(clknet_leaf_49_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload16 (.I(clknet_leaf_50_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload17 (.I(clknet_leaf_0_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload18 (.I(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload19 (.I(clknet_leaf_3_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload20 (.I(clknet_leaf_4_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 clkload21 (.I(clknet_leaf_5_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload22 (.I(clknet_leaf_6_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload23 (.I(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload24 (.I(clknet_leaf_8_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload25 (.I(clknet_leaf_9_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 clkload26 (.I(clknet_leaf_10_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 clkload27 (.I(clknet_leaf_11_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload28 (.I(clknet_leaf_47_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload29 (.I(clknet_leaf_26_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload30 (.I(clknet_leaf_27_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload31 (.I(clknet_leaf_28_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload32 (.I(clknet_leaf_29_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload33 (.I(clknet_leaf_30_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload34 (.I(clknet_leaf_32_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload35 (.I(clknet_leaf_33_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload36 (.I(clknet_leaf_34_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload37 (.I(clknet_leaf_15_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload38 (.I(clknet_leaf_16_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload39 (.I(clknet_leaf_17_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload40 (.I(clknet_leaf_18_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload41 (.I(clknet_leaf_19_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload42 (.I(clknet_leaf_21_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload43 (.I(clknet_leaf_22_clk),
    .VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_36 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_70 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_138 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_268 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_274 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_288 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_304 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_308 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_316 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_320 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_342 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_376 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_386 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_395 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_399 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_410 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_444 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_448 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_450 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_459 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_475 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_478 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_512 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_520 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_543 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_546 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_574 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_580 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_622 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_630 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_634 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_643 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_645 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_648 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_656 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_666 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_674 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_678 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_682 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_716 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_750 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_784 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_818 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_852 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_886 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_920 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_954 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_988 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_1022 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_1056 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_1090 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_1124 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_1158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_0_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_0_1226 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_0_1242 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_0_1250 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_1254 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_1_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_1_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_1_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_1_189 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_205 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_216 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_1_296 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_304 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_308 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_310 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_339 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_341 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_389 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_391 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_430 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_1_498 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_506 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_508 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_537 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_1_551 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_598 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_641 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_643 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_1_684 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_1_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_766 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_1_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_836 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_1_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_906 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_1_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_976 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_1_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_1_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_1_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_1_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_1_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_2_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_2_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_2_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_2_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_2_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_308 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_312 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_2_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_333 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_337 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_370 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_372 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_395 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_399 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_408 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_410 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_446 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_470 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_2_512 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_520 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_563 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_575 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_593 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_2_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_619 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_655 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_2_695 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_2_727 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_741 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_743 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_2_749 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_757 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_761 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_2_767 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_799 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_803 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_2_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_2_849 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_2_865 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_873 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_2_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_941 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_2_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_1011 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_2_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_2_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_2_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_2_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_2_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_2_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_3_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_3_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_3_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_162 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_164 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_3_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_3_187 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_195 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_216 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_3_235 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_267 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_269 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_288 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_3_295 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_325 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_3_336 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_344 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_348 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_3_410 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_428 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_3_439 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_447 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_3_520 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_544 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_564 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_571 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_607 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_617 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_621 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_671 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_675 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_3_681 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_697 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_699 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_714 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_718 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_720 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_726 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_728 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_741 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_754 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_3_777 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_790 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_812 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_3_821 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_829 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_870 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_880 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_884 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_908 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_3_922 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_3_954 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_3_970 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_978 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_3_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_3_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_3_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_3_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_3_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_4_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_4_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_4_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_4_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_193 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_197 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_199 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_4_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_259 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_261 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_4_273 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_281 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_4_291 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_329 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_333 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_362 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_400 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_4_410 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_424 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_438 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_4_444 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_452 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_4_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_465 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_467 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_4_510 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_518 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_522 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_4_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_561 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_590 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_608 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_646 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_650 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_4_656 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_4_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_4_683 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_780 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_4_824 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_872 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_918 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_4_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_1011 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_4_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_4_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_4_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_4_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_4_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_4_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_5_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_5_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_5_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_5_120 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_128 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_5_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_162 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_5_190 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_198 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_202 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_223 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_225 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_5_245 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_265 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_348 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_5_358 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_374 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_376 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_415 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_426 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_437 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_439 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_450 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_5_469 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_485 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_5_505 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_513 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_545 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_549 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_551 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_5_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_570 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_586 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_590 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_620 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_625 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_5_637 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_645 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_649 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_680 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_684 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_686 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_736 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_738 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_767 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_777 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_810 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_819 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_823 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_837 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_5_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_858 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_5_865 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_881 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_5_887 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_895 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_899 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_5_930 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_946 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_967 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_969 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_975 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_979 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_5_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_5_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_5_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_5_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_5_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_6_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_6_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_6_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_115 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_155 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_195 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_215 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_217 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_6_232 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_240 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_266 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_268 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_6_284 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_300 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_302 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_321 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_380 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_6_394 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_402 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_411 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_413 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_6_442 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_450 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_461 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_518 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_522 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_6_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_543 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_6_572 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_588 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_592 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_635 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_642 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_651 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_698 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_700 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_734 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_6_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_753 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_757 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_759 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_6_765 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_781 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_783 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_801 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_6_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_6_845 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_853 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_857 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_6_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_6_893 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_901 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_6_934 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_942 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_944 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_6_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_955 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_6_991 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_6_1007 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_6_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_6_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_6_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_6_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_6_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_6_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_7_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_7_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_7_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_7_120 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_128 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_132 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_147 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_165 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_175 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_214 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_7_248 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_256 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_262 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_266 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_7_290 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_306 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_7_358 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_7_394 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_410 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_483 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_485 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_501 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_7_507 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_523 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_532 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_536 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_7_552 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_7_598 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_637 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_657 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_673 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_677 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_698 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_7_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_715 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_747 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_751 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_776 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_778 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_784 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_786 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_804 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_7_811 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_819 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_835 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_848 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_873 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_907 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_909 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_7_921 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_937 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_951 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_955 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_968 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_978 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_7_994 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_7_1026 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_7_1042 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_7_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_7_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_7_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_7_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_8_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_8_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_8_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_8_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_147 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_161 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_163 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_179 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_8_188 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_204 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_231 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_259 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_309 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_313 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_321 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_8_335 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_343 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_8_373 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_8_402 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_424 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_8_442 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_450 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_8_469 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_8_485 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_510 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_512 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_8_574 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_590 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_8_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_605 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_609 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_615 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_619 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_641 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_660 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_672 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_688 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_741 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_743 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_749 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_782 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_801 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_812 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_814 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_873 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_887 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_934 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_941 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_8_974 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_8_996 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_1012 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1014 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_8_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_8_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_8_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_8_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_8_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_8_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_9_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_9_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_9_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_138 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_208 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_220 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_222 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_257 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_261 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_263 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_274 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_278 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_9_290 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_298 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_9_329 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_337 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_341 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_9_370 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_378 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_452 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_456 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_458 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_9_466 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_9_482 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_505 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_555 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_568 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_9_610 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_9_656 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_9_672 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_680 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_684 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_704 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_717 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_719 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_735 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_739 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_9_745 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_753 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_767 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_774 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_779 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_809 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_814 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_822 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_9_829 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_837 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_846 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_9_855 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_9_871 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_879 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_893 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_9_900 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_908 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_9_917 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_933 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_942 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_9_961 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_977 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_979 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_9_1006 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_9_1038 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_9_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_9_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_9_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_9_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_10_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_10_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_111 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_113 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_160 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_162 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_185 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_223 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_225 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_242 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_270 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_281 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_10_291 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_307 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_321 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_339 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_347 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_10_365 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_397 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_452 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_483 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_485 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_516 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_564 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_566 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_10_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_613 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_617 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_619 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_634 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_650 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_654 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_675 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_700 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_708 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_712 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_726 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_734 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_745 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_747 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_10_761 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_777 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_779 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_792 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_800 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_804 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_811 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_829 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_837 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_866 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_881 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_10_894 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_910 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_917 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_925 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_927 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_965 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_973 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_1012 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1014 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_10_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_10_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_10_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_10_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_10_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_10_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_11_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_11_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_11_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_112 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_11_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_208 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_226 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_230 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_11_296 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_312 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_382 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_406 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_11_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_485 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_496 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_498 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_505 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_537 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_541 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_11_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_11_596 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_11_637 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_653 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_657 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_671 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_675 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_677 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_698 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_11_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_718 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_720 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_11_738 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_802 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_806 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_11_827 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_835 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_11_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_855 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_11_873 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_881 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_883 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_11_928 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_936 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_940 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_11_970 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_978 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_11_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_11_1002 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_11_1034 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_11_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_11_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_11_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_11_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_12_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_12_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_12_69 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_12_85 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_93 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_97 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_111 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_12_151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_159 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_12_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_185 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_249 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_312 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_340 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_361 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_12_393 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_409 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_12_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_469 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_490 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_531 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_588 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_592 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_12_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_605 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_607 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_626 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_630 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_646 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_650 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_652 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_685 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_694 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_707 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_711 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_713 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_734 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_12_742 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_750 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_12_758 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_12_774 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_782 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_803 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_12_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_815 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_12_838 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_846 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_850 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_852 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_12_865 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_873 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_881 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_883 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_903 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_12_930 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_938 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_942 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_944 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_951 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_12_968 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_12_984 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_997 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1014 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_12_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_12_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_12_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_12_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_12_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_12_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_13_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_13_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_13_124 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_132 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_13_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_13_166 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_178 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_13_189 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_197 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_207 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_13_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_220 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_224 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_226 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_240 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_273 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_277 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_13_302 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_310 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_13_334 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_356 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_358 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_385 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_455 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_465 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_469 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_478 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_482 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_13_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_13_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_540 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_544 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_557 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_564 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_627 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_13_655 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_691 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_693 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_13_710 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_718 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_722 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_13_746 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_754 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_13_777 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_793 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_795 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_801 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_813 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_817 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_838 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_13_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_13_875 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_883 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_905 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_909 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_13_917 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_942 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_13_954 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_962 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_990 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_992 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_13_1021 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_13_1037 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_1045 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_1049 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_13_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_13_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_13_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_13_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_14_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_14_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_14_127 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_143 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_14_155 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_163 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_167 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_169 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_199 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_14_215 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_223 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_229 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_238 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_257 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_14_286 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_14_302 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_14_325 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_341 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_14_404 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_436 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_14_462 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_470 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_474 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_491 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_14_505 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_539 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_14_549 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_557 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_561 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_572 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_576 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_14_641 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_14_657 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_682 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_686 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_688 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_14_712 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_720 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_14_743 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_780 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_784 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_881 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_14_890 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_911 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_915 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_957 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_961 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_963 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_968 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_984 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_988 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_990 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_1009 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_1013 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_14_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_1025 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_14_1059 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_14_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_14_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_14_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_14_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_14_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_15_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_15_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_92 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_94 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_99 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_131 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_165 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_189 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_15_197 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_205 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_220 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_224 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_15_238 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_15_254 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_262 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_266 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_268 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_277 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_15_287 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_323 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_339 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_354 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_365 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_405 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_407 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_417 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_428 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_430 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_463 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_15_509 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_517 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_557 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_15_647 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_679 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_696 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_15_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_710 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_15_719 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_727 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_731 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_15_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_745 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_15_778 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_786 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_790 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_812 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_816 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_818 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_824 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_826 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_15_850 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_866 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_870 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_893 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_897 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_908 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_15_922 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_943 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_945 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_15_958 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_974 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_978 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_991 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_995 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_997 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_15_1012 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_1044 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_1048 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_15_1108 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_15_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_15_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_15_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_16_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_16_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_53 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_16_124 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_140 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_144 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_152 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_156 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_16_167 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_16_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_193 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_195 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_218 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_231 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_267 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_16_291 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_307 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_309 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_348 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_374 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_395 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_428 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_430 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_16_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_465 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_16_474 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_16_498 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_16_514 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_522 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_16_544 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_552 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_16_577 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_593 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_16_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_605 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_607 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_16_623 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_639 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_16_654 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_662 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_701 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_703 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_732 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_734 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_16_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_753 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_757 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_16_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_804 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_16_867 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_16_928 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_944 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_16_957 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_965 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_974 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_978 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_16_1005 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1013 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_16_1047 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_1055 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_1059 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1061 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_16_1072 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_1080 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1084 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_16_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_16_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_16_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_16_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_16_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_17_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_83 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_17_93 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_17_124 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_17_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_17_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_217 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_263 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_267 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_17_295 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_303 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_340 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_344 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_364 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_368 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_398 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_402 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_17_435 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_443 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_447 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_449 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_17_504 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_520 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_17_542 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_558 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_566 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_580 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_584 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_17_590 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_598 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_628 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_17_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_640 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_644 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_646 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_688 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_692 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_699 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_17_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_710 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_17_716 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_745 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_749 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_751 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_17_757 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_765 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_777 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_779 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_835 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_17_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_850 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_852 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_909 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_17_917 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_925 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_929 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_931 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_944 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_946 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_954 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_975 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_979 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_17_1013 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_1029 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_17_1042 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_17_1082 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_1114 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_1118 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_17_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_17_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_17_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_18_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_18_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_53 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_57 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_115 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_146 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_18_199 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_215 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_219 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_224 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_233 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_235 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_242 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_18_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_18_263 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_271 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_275 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_295 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_304 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_306 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_18_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_333 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_356 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_18_370 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_378 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_382 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_18_393 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_18_425 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_18_441 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_449 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_453 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_480 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_482 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_18_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_570 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_18_603 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_619 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_623 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_625 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_18_656 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_715 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_717 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_761 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_815 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_18_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_885 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_889 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_909 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_923 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_944 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_959 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_963 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_18_977 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_985 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_989 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_18_1006 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1014 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_1047 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_18_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_18_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_18_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_18_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_18_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_19_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_19_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_50 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_74 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_103 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_137 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_149 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_160 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_233 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_19_240 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_248 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_19_260 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_268 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_270 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_277 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_290 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_361 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_19_377 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_19_393 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_401 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_416 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_19_430 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_438 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_442 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_456 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_460 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_488 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_505 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_507 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_520 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_557 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_19_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_570 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_584 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_588 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_590 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_19_609 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_625 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_691 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_731 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_735 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_749 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_753 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_19_759 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_767 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_19_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_785 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_837 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_19_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_19_882 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_898 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_900 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_906 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_914 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_19_920 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_928 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_932 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_19_938 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_946 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_948 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_19_957 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_973 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_977 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_979 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_19_1004 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_1012 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_19_1039 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1047 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1049 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1056 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_19_1093 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_19_1109 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_1117 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_1119 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_19_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_19_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_19_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_20_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_20_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_20_69 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_77 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_91 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_95 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_103 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_20_120 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_128 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_132 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_20_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_173 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_239 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_249 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_280 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_350 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_424 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_453 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_461 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_503 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_507 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_514 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_522 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_531 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_533 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_20_552 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_560 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_610 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_20_641 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_20_722 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_730 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_734 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_745 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_747 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_20_768 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_776 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_783 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_790 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_802 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_804 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_838 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_844 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_860 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_20_918 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_926 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_930 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_943 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_953 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_955 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_962 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_20_972 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_980 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_20_1002 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_1010 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1014 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_20_1039 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_1047 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1051 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1053 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1083 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_20_1109 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_20_1141 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_1149 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_1153 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_20_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_20_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_20_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_20_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_21_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_21_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_106 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_21_114 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_126 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_137 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_21_155 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_230 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_298 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_343 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_21_386 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_394 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_396 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_21_434 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_442 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_21_473 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_500 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_502 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_515 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_532 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_21_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_570 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_574 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_576 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_595 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_599 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_608 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_675 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_679 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_690 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_692 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_711 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_715 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_740 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_744 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_21_780 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_796 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_21_824 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_21_872 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_21_888 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_896 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_898 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_904 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_908 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_916 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_918 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_949 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_951 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_976 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_986 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_21_1000 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1008 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1010 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_21_1035 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_1043 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1047 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1049 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_21_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_1068 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_21_1073 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_1089 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_21_1112 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_21_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_21_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_21_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_22_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_22_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_53 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_55 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_84 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_121 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_22_164 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_182 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_22_190 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_198 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_205 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_207 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_222 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_224 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_273 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_275 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_347 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_351 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_353 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_383 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_22_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_22_424 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_22_440 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_448 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_452 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_461 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_463 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_482 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_22_498 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_514 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_516 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_22_539 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_22_555 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_563 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_567 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_22_576 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_592 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_646 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_662 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_672 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_676 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_678 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_22_696 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_22_712 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_720 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_724 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_726 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_733 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_22_742 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_750 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_754 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_22_766 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_799 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_803 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_809 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_815 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_817 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_838 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_850 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_22_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_885 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_889 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_22_914 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_930 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_943 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_952 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_956 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_22_980 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_996 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1000 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1037 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1064 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1074 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1076 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_22_1101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_22_1133 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_1149 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_1153 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_22_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_22_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_22_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_22_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_23_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_96 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_152 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_160 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_164 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_199 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_207 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_277 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_287 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_338 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_354 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_390 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_394 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_23_430 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_487 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_508 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_515 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_523 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_552 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_570 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_595 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_599 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_601 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_608 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_627 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_640 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_657 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_683 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_689 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_697 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_699 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_707 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_23_725 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_757 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_765 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_774 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_813 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_847 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_855 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_880 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_884 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_886 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_23_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_928 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_936 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_946 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_954 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_963 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_967 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_979 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_23_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_990 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_998 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_1035 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_23_1104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_23_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_23_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_23_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_24_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_24_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_24_69 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_77 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_93 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_97 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_24_123 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_24_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_191 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_220 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_253 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_326 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_379 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_383 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_392 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_453 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_462 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_508 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_512 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_24_547 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_563 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_615 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_619 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_621 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_24_630 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_700 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_732 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_734 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_776 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_798 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_802 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_804 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_24_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_815 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_24_836 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_852 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_870 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_24_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_931 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_24_971 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_1003 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1007 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1013 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1044 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1060 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1062 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_24_1076 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1084 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_24_1098 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_24_1130 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_24_1146 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1154 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_24_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_24_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_24_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_24_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_25_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_25_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_92 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_105 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_114 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_118 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_137 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_146 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_148 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_25_196 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_204 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_208 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_258 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_260 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_269 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_271 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_347 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_25_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_388 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_397 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_417 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_25_428 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_436 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_440 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_488 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_25_500 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_528 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_25_534 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_542 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_556 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_585 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_589 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_25_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_648 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_650 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_670 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_724 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_726 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_755 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_759 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_765 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_25_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_788 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_795 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_799 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_25_809 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_25_825 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_833 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_837 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_846 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_850 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_25_871 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_25_887 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_895 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_909 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_25_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_928 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_951 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_964 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_974 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_978 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_25_1012 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_1020 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1024 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1038 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1049 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_25_1057 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1065 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_25_1073 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_1089 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_25_1103 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_1119 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_25_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_25_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_25_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_26_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_26_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_53 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_168 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_185 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_205 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_211 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_252 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_260 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_286 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_292 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_294 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_313 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_326 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_334 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_336 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_353 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_355 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_26_364 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_405 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_432 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_440 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_448 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_452 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_461 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_491 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_533 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_26_570 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_586 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_623 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_631 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_675 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_679 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_681 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_715 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_723 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_26_765 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_781 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_802 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_804 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_819 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_831 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_833 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_864 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_872 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_885 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_917 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_925 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_934 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_943 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_953 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_957 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_26_966 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_26_998 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1014 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_1029 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1033 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1035 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_1048 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_1056 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_1080 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1084 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_26_1113 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_1145 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_1153 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_26_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_26_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_26_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_26_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_27_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_27_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_27_50 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_58 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_62 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_64 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_138 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_27_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_154 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_27_184 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_27_200 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_208 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_220 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_27_225 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_233 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_235 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_248 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_252 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_268 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_272 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_274 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_290 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_27_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_322 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_417 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_459 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_487 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_27_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_528 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_530 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_543 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_545 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_27_550 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_558 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_27_585 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_593 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_595 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_628 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_27_662 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_670 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_27_710 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_718 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_732 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_751 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_755 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_757 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_776 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_818 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_834 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_838 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_855 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_859 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_861 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_866 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_876 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_893 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_897 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_935 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_27_952 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_27_968 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_976 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_27_1012 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1020 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1057 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1059 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1077 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1079 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1100 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_27_1109 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_1117 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_1119 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_27_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_27_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_27_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_28_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_28_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_69 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_73 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_149 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_193 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_195 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_28_252 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_260 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_262 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_28_300 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_308 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_312 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_28_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_330 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_348 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_28_365 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_28_405 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_28_421 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_429 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_448 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_452 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_471 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_473 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_28_485 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_28_501 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_509 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_552 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_554 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_560 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_564 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_602 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_622 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_28_654 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_662 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_28_677 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_693 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_28_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_718 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_722 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_729 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_733 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_28_760 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_776 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_778 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_28_794 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_802 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_804 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_28_813 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_845 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_855 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_859 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_861 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_889 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_893 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_917 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_931 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_28_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_963 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1013 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1034 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_28_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1054 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_28_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_1148 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_1152 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1154 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_28_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_28_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_28_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_28_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_29_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_76 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_159 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_207 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_29_259 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_267 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_271 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_29_298 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_306 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_326 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_29_392 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_400 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_404 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_459 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_29_500 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_508 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_510 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_587 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_608 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_612 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_625 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_29_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_648 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_652 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_654 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_29_691 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_699 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_29_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_710 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_712 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_29_760 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_768 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_776 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_806 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_29_820 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_828 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_830 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_866 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_875 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_906 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_29_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_928 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_932 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_29_961 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_969 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_973 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_29_1037 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_1045 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1049 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_29_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_29_1084 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_1092 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_1096 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1098 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_29_1111 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_1119 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_29_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_29_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_29_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_30_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_30_67 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_75 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_77 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_30_88 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_30_165 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_173 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_30_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_30_193 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_201 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_205 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_30_228 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_30_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_257 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_283 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_285 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_294 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_308 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_30_325 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_357 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_361 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_371 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_412 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_30_439 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_520 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_529 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_592 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_30_613 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_30_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_671 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_703 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_705 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_715 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_724 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_726 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_732 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_734 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_744 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_746 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_764 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_768 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_784 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_803 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_30_821 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_841 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_845 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_847 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_856 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_860 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_862 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_871 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_30_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_30_917 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_30_933 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_941 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_30_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_963 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1000 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1002 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1035 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1041 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1056 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1058 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_1071 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1075 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1093 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1095 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_30_1100 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_30_1132 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_1148 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_1152 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1154 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_30_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_30_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_30_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_30_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_31_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_38 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_40 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_51 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_59 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_69 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_80 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_31_112 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_128 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_132 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_134 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_155 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_163 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_197 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_205 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_31_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_228 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_236 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_249 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_257 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_267 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_271 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_301 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_309 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_324 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_332 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_414 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_446 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_458 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_467 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_475 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_477 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_500 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_538 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_540 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_553 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_557 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_598 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_658 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_662 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_694 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_698 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_717 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_719 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_735 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_749 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_757 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_795 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_797 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_815 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_819 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_832 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_850 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_854 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_856 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_909 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_927 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_935 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_966 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1000 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1002 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_1036 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_31_1105 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_1113 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_1117 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_1119 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_31_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_31_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_31_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_30 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_32_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_45 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_32_76 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_96 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_32_117 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_125 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_129 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_32_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_32_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_32_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_185 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_189 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_259 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_269 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_325 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_329 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_379 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_383 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_32_403 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_446 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_32_478 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_494 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_535 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_537 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_32_550 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_558 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_564 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_32_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_32_613 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_621 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_623 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_32_652 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_660 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_32_683 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_699 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_703 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_732 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_734 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_742 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_794 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_798 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_815 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_819 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_821 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_826 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_32_854 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_862 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_872 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_32_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_885 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_887 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_32_894 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_902 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_906 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_908 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_931 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_32_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_963 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_967 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_969 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_1009 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1013 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1042 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_32_1062 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_1078 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1082 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1084 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_32_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_1148 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_1152 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1154 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_32_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_32_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_32_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_32_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_10 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_33_46 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_62 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_68 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_76 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_78 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_110 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_146 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_159 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_161 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_33_190 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_220 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_256 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_260 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_301 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_328 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_344 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_348 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_369 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_377 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_383 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_395 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_33_432 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_485 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_500 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_525 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_558 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_33_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_578 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_586 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_588 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_617 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_625 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_636 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_638 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_648 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_662 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_670 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_672 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_687 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_691 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_693 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_712 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_726 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_730 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_760 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_816 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_824 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_850 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_871 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_873 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_886 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_898 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_902 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_904 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_957 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_965 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_969 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_1000 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_33_1031 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1047 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1049 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_1060 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1064 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_33_1075 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1091 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_1093 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_33_1106 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_1114 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_1118 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_33_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_33_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_33_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_32 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_55 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_57 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_80 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_102 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_148 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_179 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_34_208 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_224 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_233 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_261 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_289 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_293 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_306 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_34_325 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_333 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_337 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_371 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_405 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_407 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_413 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_417 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_426 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_428 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_34_433 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_449 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_453 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_494 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_496 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_34_578 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_34_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_34_617 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_625 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_657 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_659 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_727 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_739 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_794 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_798 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_800 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_821 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_823 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_34_828 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_836 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_840 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_34_862 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_887 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_891 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_34_904 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_944 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_979 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1000 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1002 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_34_1029 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_1037 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_1071 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1075 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1084 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1089 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_34_1110 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_34_1142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_1150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1154 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_34_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_34_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_34_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_34_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_35_55 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_59 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_61 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_35_85 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_93 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_95 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_124 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_35_133 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_137 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_35_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_35_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_154 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_190 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_204 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_35_316 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_324 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_35_331 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_35_339 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_343 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_354 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_376 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_383 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_35_404 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_412 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_35_440 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_35_472 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_488 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_35_572 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_35_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_35_640 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_644 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_35_652 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_660 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_698 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_35_732 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_740 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_35_750 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_758 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_35_785 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_789 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_804 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_35_831 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_844 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_858 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_860 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_35_905 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_909 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_914 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_920 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_927 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_1030 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_1032 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_35_1088 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_35_1100 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_35_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_35_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_35_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_35_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_36_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_18 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_31 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_36_45 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_53 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_36_83 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_109 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_36_118 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_126 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_130 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_36_159 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_183 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_203 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_207 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_36_213 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_225 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_242 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_249 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_296 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_307 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_309 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_36_337 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_345 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_382 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_36_399 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_459 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_36_466 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_482 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_523 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_529 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_558 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_592 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_36_622 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_638 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_640 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_36_649 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_662 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_700 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_36_727 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_36_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_753 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_36_793 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_801 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_36_821 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_829 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_833 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_36_855 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_871 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_904 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_908 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_940 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_944 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_36_967 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_983 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_1005 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1009 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_36_1023 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_1031 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1043 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1049 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_1058 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1074 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1082 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1084 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_36_1097 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_36_1129 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_36_1145 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_1153 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_36_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_36_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_36_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_36_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_56 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_82 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_86 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_37_96 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_108 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_113 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_124 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_128 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_156 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_37_164 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_180 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_182 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_205 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_218 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_220 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_231 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_272 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_305 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_37_329 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_337 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_341 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_358 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_37_389 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_405 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_407 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_424 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_37_439 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_37_576 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_584 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_588 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_590 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_607 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_611 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_613 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_636 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_657 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_37_722 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_738 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_757 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_37_795 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_803 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_37_829 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_837 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_37_852 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_860 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_862 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_880 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_884 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_886 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_37_899 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_907 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_909 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_37_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_920 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_922 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_932 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_951 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_37_994 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_1025 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1039 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1074 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_37_1099 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_1115 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_1119 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_37_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_37_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_37_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_38_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_10 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_14 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_16 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_48 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_52 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_103 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_156 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_38_323 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_331 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_335 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_337 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_358 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_373 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_398 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_402 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_421 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_430 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_465 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_479 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_483 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_522 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_544 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_38_584 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_592 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_38_643 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_659 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_685 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_687 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_719 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_728 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_732 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_734 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_38_749 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_757 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_767 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_771 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_38_791 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_799 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_803 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_821 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_38_835 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_851 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_855 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_868 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_872 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_38_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_38_893 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_901 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_905 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_919 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_958 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_38_989 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_997 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1001 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_38_1064 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_1080 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1084 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_38_1092 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_38_1124 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_38_1140 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_1148 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_1152 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1154 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_38_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_38_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_38_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_38_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_39_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_39_38 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_76 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_93 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_164 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_166 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_185 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_195 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_208 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_231 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_242 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_278 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_298 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_302 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_327 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_329 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_39_339 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_347 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_39_360 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_368 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_378 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_380 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_391 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_39_428 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_436 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_39_444 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_471 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_473 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_499 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_536 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_571 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_573 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_39_593 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_601 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_610 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_39_617 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_625 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_39_640 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_648 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_650 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_39_684 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_39_710 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_718 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_722 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_39_756 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_764 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_768 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_776 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_799 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_810 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_812 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_821 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_39_831 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_867 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_869 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_878 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_880 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_904 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_908 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_925 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_939 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_941 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_950 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_39_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_39_1027 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_1043 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_1047 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_1049 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_39_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_39_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_39_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_39_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_40_49 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_57 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_74 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_76 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_99 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_103 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_160 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_173 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_40_207 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_239 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_40_292 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_300 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_321 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_342 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_348 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_40_377 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_402 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_470 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_474 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_40_490 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_40_506 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_40_583 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_609 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_611 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_653 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_40_675 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_691 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_40_720 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_728 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_732 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_734 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_752 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_771 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_802 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_804 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_40_815 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_851 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_40_858 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_40_909 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_917 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_926 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_928 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_939 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_943 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_952 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_964 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_40_998 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1014 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_40_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_40_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_40_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_40_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_40_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_40_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_41_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_18 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_41_43 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_51 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_55 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_87 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_130 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_160 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_226 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_41_235 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_245 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_276 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_286 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_301 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_324 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_328 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_41_337 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_345 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_41_386 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_402 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_413 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_417 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_41_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_453 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_455 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_41_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_500 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_504 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_523 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_549 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_577 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_617 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_658 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_675 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_693 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_699 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_41_714 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_41_758 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_766 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_41_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_780 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_782 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_41_800 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_816 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_850 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_881 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_41_887 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_903 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_907 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_909 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_918 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_942 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_41_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_41_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_41_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_41_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_41_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_42_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_18 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_22 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_24 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_33 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_42_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_45 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_67 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_71 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_42_91 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_99 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_103 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_111 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_113 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_124 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_153 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_42_219 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_239 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_259 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_42_271 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_308 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_312 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_42_331 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_347 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_359 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_363 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_42_377 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_396 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_400 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_42_431 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_452 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_42_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_465 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_42_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_497 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_42_573 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_589 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_593 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_42_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_613 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_617 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_654 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_656 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_690 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_42_750 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_42_782 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_798 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_802 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_804 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_42_816 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_832 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_834 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_42_840 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_856 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_858 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_868 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_872 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_42_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_885 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_891 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_42_904 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_949 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_42_978 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_1010 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1014 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_42_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_42_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_42_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_42_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_42_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_42_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_43_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_10 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_14 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_43_49 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_57 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_85 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_137 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_180 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_204 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_208 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_43_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_220 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_248 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_252 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_262 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_264 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_273 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_277 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_43_292 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_300 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_340 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_342 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_360 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_43_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_389 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_436 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_43_472 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_488 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_43_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_573 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_603 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_605 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_43_649 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_657 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_690 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_694 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_704 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_43_713 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_729 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_731 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_752 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_756 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_777 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_798 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_823 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_43_854 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_870 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_43_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_920 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_922 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_931 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_43_960 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_976 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_43_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_43_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_43_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_43_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_43_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_123 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_162 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_223 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_239 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_261 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_263 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_44_294 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_302 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_306 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_347 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_44_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_454 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_520 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_561 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_44_575 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_625 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_44_636 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_44_652 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_660 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_674 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_44_688 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_696 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_700 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_44_706 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_719 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_723 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_729 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_44_762 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_770 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_801 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_44_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_856 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_871 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_890 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_44_924 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_940 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_944 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_44_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_1011 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_44_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_44_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_44_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_44_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_44_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_44_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_45_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_30 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_32 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_43 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_51 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_68 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_82 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_95 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_130 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_201 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_220 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_224 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_246 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_257 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_261 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_263 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_278 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_45_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_298 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_318 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_320 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_358 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_388 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_396 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_400 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_402 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_428 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_468 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_510 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_518 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_537 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_545 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_549 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_558 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_45_578 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_621 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_45_653 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_697 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_699 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_707 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_718 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_729 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_757 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_765 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_780 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_45_795 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_811 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_820 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_829 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_837 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_850 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_897 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_905 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_909 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_45_918 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_45_950 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_45_966 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_974 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_978 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_45_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_45_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_45_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_45_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_45_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_46_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_18 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_22 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_53 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_61 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_63 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_94 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_102 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_127 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_135 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_213 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_217 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_249 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_286 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_294 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_298 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_306 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_46_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_333 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_46_354 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_382 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_397 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_405 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_417 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_431 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_439 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_453 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_46_474 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_46_506 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_522 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_529 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_46_535 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_551 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_555 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_557 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_586 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_621 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_625 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_627 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_661 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_671 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_686 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_693 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_701 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_705 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_730 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_734 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_46_760 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_776 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_780 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_782 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_788 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_835 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_843 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_847 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_860 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_868 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_872 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_879 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_887 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_895 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_899 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_46_924 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_940 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_944 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_46_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_1011 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_46_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_46_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_46_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_46_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_46_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_46_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_59 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_67 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_69 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_47_95 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_111 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_127 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_135 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_144 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_161 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_168 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_176 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_216 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_347 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_375 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_385 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_393 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_397 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_410 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_439 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_447 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_481 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_506 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_512 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_531 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_570 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_580 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_584 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_599 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_603 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_605 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_616 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_624 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_628 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_634 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_47_656 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_672 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_680 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_687 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_696 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_711 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_47_720 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_752 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_760 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_812 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_816 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_822 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_830 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_834 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_859 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_863 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_887 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_895 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_899 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_909 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_47_919 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_47_951 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_47_967 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_975 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_979 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_47_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_47_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_47_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_47_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_47_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_48_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_18 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_22 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_54 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_62 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_76 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_84 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_92 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_100 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_193 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_201 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_205 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_215 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_223 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_229 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_236 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_238 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_249 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_298 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_302 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_309 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_313 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_321 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_339 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_343 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_375 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_383 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_395 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_397 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_425 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_433 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_463 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_469 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_546 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_554 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_579 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_583 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_592 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_627 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_635 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_652 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_660 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_675 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_710 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_714 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_716 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_729 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_733 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_745 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_763 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_765 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_774 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_785 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_804 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_809 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_827 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_831 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_833 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_858 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_862 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_864 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_885 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_889 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_48_925 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_941 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_48_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_1011 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_48_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_48_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_48_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_48_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_48_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_48_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_49_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_18 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_49_50 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_86 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_105 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_115 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_49_122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_138 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_49_183 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_203 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_222 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_49_239 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_286 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_288 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_49_334 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_354 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_361 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_49_383 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_399 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_426 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_436 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_522 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_49_546 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_554 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_558 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_570 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_572 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_49_579 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_595 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_599 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_628 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_636 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_666 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_694 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_698 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_706 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_49_720 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_728 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_732 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_49_759 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_767 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_804 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_806 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_49_831 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_49_857 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_873 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_880 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_49_889 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_49_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_976 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_49_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_49_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_49_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_49_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_49_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_30 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_55 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_59 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_50_87 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_103 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_50_119 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_50_135 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_143 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_153 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_50_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_205 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_224 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_298 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_50_322 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_50_338 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_346 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_350 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_382 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_384 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_50_392 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_400 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_417 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_436 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_451 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_475 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_479 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_481 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_510 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_520 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_50_552 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_560 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_564 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_566 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_50_578 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_640 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_50_651 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_659 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_663 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_733 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_739 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_50_752 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_768 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_774 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_50_784 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_800 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_804 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_50_816 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_50_832 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_868 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_872 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_893 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_50_907 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_939 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_943 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_50_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_1011 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_50_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_50_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_50_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_50_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_50_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_50_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_51_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_51_10 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_14 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_67 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_69 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_51_94 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_51_128 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_51_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_51_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_160 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_51_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_51_180 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_184 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_204 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_51_221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_51_243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_277 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_51_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_286 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_288 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_315 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_348 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_388 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_390 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_403 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_405 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_446 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_51_481 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_505 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_507 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_554 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_51_586 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_629 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_655 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_697 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_699 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_51_724 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_51_761 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_794 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_51_823 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_831 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_839 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_850 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_852 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_51_861 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_51_886 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_51_902 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_51_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_51_976 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_51_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_51_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_51_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_51_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_51_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_51_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_51_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_10 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_14 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_32 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_55 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_59 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_94 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_102 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_109 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_127 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_143 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_181 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_189 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_193 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_52_215 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_231 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_239 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_311 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_356 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_358 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_393 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_413 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_449 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_453 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_482 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_490 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_498 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_502 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_504 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_513 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_535 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_539 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_541 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_52_547 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_563 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_593 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_630 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_638 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_642 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_660 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_52_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_683 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_689 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_699 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_713 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_726 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_734 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_753 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_761 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_763 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_780 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_797 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_52_817 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_833 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_841 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_843 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_52_850 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_866 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_874 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_52_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_941 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_52_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_1011 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_52_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_52_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_52_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_52_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_52_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_52_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_53_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_18 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_22 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_24 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_53_35 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_53_51 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_103 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_53_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_150 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_175 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_53_194 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_53_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_220 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_296 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_300 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_53_329 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_345 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_53_379 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_53_412 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_53_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_53_438 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_446 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_450 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_53_460 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_476 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_480 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_53_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_500 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_502 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_53_526 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_554 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_558 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_53_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_570 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_53_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_648 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_652 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_53_681 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_697 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_699 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_53_707 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_53_739 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_53_755 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_763 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_767 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_769 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_778 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_53_790 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_53_822 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_838 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_53_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_906 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_53_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_976 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_53_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_53_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_53_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_53_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_53_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_54_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_68 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_54_93 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_111 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_54_135 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_143 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_173 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_205 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_242 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_253 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_298 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_302 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_317 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_54_330 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_338 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_340 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_357 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_361 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_371 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_54_377 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_54_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_395 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_54_410 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_429 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_431 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_479 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_481 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_521 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_529 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_54_563 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_571 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_575 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_591 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_54_603 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_611 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_615 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_617 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_54_646 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_662 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_54_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_731 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_54_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_801 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_54_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_871 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_54_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_941 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_54_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_1011 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_54_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_54_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_54_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_54_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_54_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_54_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_55_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_55_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_80 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_82 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_55_87 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_95 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_97 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_55_126 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_134 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_138 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_55_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_176 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_178 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_197 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_199 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_216 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_258 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_55_267 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_275 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_279 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_55_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_298 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_302 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_304 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_327 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_343 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_347 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_55_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_360 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_55_383 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_431 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_435 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_448 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_55_461 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_469 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_479 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_489 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_55_492 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_500 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_520 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_55_529 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_545 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_558 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_55_618 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_626 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_55_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_696 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_55_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_766 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_55_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_836 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_55_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_906 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_55_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_976 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_55_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_55_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_55_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_55_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_55_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_56_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_56_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_56_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_56_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_147 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_149 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_56_160 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_168 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_205 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_56_215 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_223 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_229 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_240 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_56_273 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_281 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_56_297 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_313 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_329 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_333 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_368 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_381 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_391 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_56_413 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_56_437 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_445 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_465 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_467 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_499 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_503 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_56_580 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_588 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_592 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_56_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_605 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_609 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_611 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_56_640 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_56_656 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_56_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_731 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_56_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_801 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_56_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_871 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_56_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_941 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_56_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_1011 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_56_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_56_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_56_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_56_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_56_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_56_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_57_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_57_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_57_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_57_174 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_182 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_57_189 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_205 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_209 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_268 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_284 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_57_315 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_323 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_327 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_329 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_360 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_362 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_57_385 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_393 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_414 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_418 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_57_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_430 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_446 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_450 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_57_464 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_472 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_476 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_57_497 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_513 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_517 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_57_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_535 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_57_545 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_553 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_557 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_57_570 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_624 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_628 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_57_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_696 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_57_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_766 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_57_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_836 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_57_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_906 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_57_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_976 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_57_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_57_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_57_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_57_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_57_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_58_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_58_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_58_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_171 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_58_177 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_241 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_58_247 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_58_263 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_271 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_58_307 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_343 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_349 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_365 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_58_375 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_383 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_58_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_395 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_397 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_58_421 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_429 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_431 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_58_465 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_473 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_503 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_517 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_519 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_527 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_529 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_542 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_58_558 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_590 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_594 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_601 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_58_628 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_660 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_664 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_58_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_731 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_58_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_801 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_58_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_871 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_58_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_941 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_58_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_1011 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_58_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_58_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_58_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_58_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_58_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_58_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_59_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_66 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_59_72 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_136 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_59_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_59_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_59_244 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_252 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_59_262 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_278 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_59_282 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_344 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_348 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_59_352 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_360 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_362 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_419 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_422 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_444 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_469 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_473 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_59_549 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_557 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_559 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_59_562 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_626 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_59_632 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_696 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_59_702 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_766 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_59_772 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_836 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_59_842 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_906 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_59_912 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_976 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_59_982 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_1046 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_59_1052 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_1116 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_59_1122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_59_1186 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_59_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_60_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_34 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_60_37 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_101 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_60_107 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_60_139 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_60_155 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_163 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_173 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_185 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_189 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_199 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_203 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_212 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_216 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_225 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_277 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_281 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_312 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_314 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_323 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_357 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_361 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_387 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_457 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_60_466 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_482 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_486 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_508 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_518 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_522 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_524 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_539 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_543 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_60_573 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_589 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_593 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_60_597 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_661 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_60_667 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_731 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_60_737 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_801 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_60_807 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_871 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_60_877 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_941 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_60_947 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_1011 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_60_1017 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_1081 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_60_1087 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_1151 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_64 FILLER_60_1157 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_1221 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_60_1227 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_60_1243 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_60_1251 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_1255 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_2 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_61_36 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_52 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_61_57 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_65 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_67 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_61_74 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_78 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_61_83 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_91 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_61_96 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_100 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_104 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_61_109 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_117 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_61_122 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_130 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_135 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_61_138 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_142 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_61_148 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_61_164 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_168 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_172 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_206 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_240 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_304 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_338 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_342 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_61_376 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_392 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_61_398 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_406 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_410 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_444 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_478 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_512 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_546 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_61_600 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_61_608 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_614 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_648 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_682 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_716 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_750 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_784 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_818 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_852 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_886 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_920 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_954 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_988 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_1022 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_1056 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_1090 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_1124 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_1158 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_32 FILLER_61_1192 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_16 FILLER_61_1226 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_8 FILLER_61_1242 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fillcap_4 FILLER_61_1250 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_1254 (.VDD(VPWR),
    .VNW(VPWR),
    .VPW(VGND),
    .VSS(VGND));
 assign uio_oe[0] = net173;
 assign uio_oe[1] = net174;
 assign uio_oe[2] = net175;
 assign uio_oe[3] = net176;
 assign uio_oe[4] = net177;
 assign uio_oe[5] = net178;
 assign uio_oe[6] = net179;
 assign uio_oe[7] = net180;
endmodule
